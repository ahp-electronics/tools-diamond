library verilog;
use verilog.vl_types.all;
entity ESBA is
    generic(
        UDS_TRN         : string  := "LSCC_UDS_TRN_VAL";
        UDS_TRN_FORMAT  : string  := "ASCII"
    );
    port(
        WBDATO31        : out    vl_logic;
        WBDATO30        : out    vl_logic;
        WBDATO29        : out    vl_logic;
        WBDATO28        : out    vl_logic;
        WBDATO27        : out    vl_logic;
        WBDATO26        : out    vl_logic;
        WBDATO25        : out    vl_logic;
        WBDATO24        : out    vl_logic;
        WBDATO23        : out    vl_logic;
        WBDATO22        : out    vl_logic;
        WBDATO21        : out    vl_logic;
        WBDATO20        : out    vl_logic;
        WBDATO19        : out    vl_logic;
        WBDATO18        : out    vl_logic;
        WBDATO17        : out    vl_logic;
        WBDATO16        : out    vl_logic;
        WBDATO15        : out    vl_logic;
        WBDATO14        : out    vl_logic;
        WBDATO13        : out    vl_logic;
        WBDATO12        : out    vl_logic;
        WBDATO11        : out    vl_logic;
        WBDATO10        : out    vl_logic;
        WBDATO9         : out    vl_logic;
        WBDATO8         : out    vl_logic;
        WBDATO7         : out    vl_logic;
        WBDATO6         : out    vl_logic;
        WBDATO5         : out    vl_logic;
        WBDATO4         : out    vl_logic;
        WBDATO3         : out    vl_logic;
        WBDATO2         : out    vl_logic;
        WBDATO1         : out    vl_logic;
        WBDATO0         : out    vl_logic;
        WBDATI31        : in     vl_logic;
        WBDATI30        : in     vl_logic;
        WBDATI29        : in     vl_logic;
        WBDATI28        : in     vl_logic;
        WBDATI27        : in     vl_logic;
        WBDATI26        : in     vl_logic;
        WBDATI25        : in     vl_logic;
        WBDATI24        : in     vl_logic;
        WBDATI23        : in     vl_logic;
        WBDATI22        : in     vl_logic;
        WBDATI21        : in     vl_logic;
        WBDATI20        : in     vl_logic;
        WBDATI19        : in     vl_logic;
        WBDATI18        : in     vl_logic;
        WBDATI17        : in     vl_logic;
        WBDATI16        : in     vl_logic;
        WBDATI15        : in     vl_logic;
        WBDATI14        : in     vl_logic;
        WBDATI13        : in     vl_logic;
        WBDATI12        : in     vl_logic;
        WBDATI11        : in     vl_logic;
        WBDATI10        : in     vl_logic;
        WBDATI9         : in     vl_logic;
        WBDATI8         : in     vl_logic;
        WBDATI7         : in     vl_logic;
        WBDATI6         : in     vl_logic;
        WBDATI5         : in     vl_logic;
        WBDATI4         : in     vl_logic;
        WBDATI3         : in     vl_logic;
        WBDATI2         : in     vl_logic;
        WBDATI1         : in     vl_logic;
        WBDATI0         : in     vl_logic;
        WBSTBI          : in     vl_logic;
        WBCLKI          : in     vl_logic;
        ASFCLKI         : in     vl_logic;
        WBRSTI          : in     vl_logic;
        ASFRESETI       : in     vl_logic;
        WBADRI17        : in     vl_logic;
        WBADRI16        : in     vl_logic;
        WBADRI15        : in     vl_logic;
        WBADRI14        : in     vl_logic;
        WBADRI13        : in     vl_logic;
        WBADRI12        : in     vl_logic;
        WBADRI11        : in     vl_logic;
        WBADRI10        : in     vl_logic;
        WBADRI9         : in     vl_logic;
        WBADRI8         : in     vl_logic;
        WBADRI7         : in     vl_logic;
        WBADRI6         : in     vl_logic;
        WBADRI5         : in     vl_logic;
        WBADRI4         : in     vl_logic;
        WBADRI3         : in     vl_logic;
        WBADRI2         : in     vl_logic;
        WBADRI1         : in     vl_logic;
        WBADRI0         : in     vl_logic;
        WBACKO          : out    vl_logic;
        ASFFULLO        : out    vl_logic;
        ASFEMPTYO       : out    vl_logic;
        WBCYCI          : in     vl_logic;
        WBWEI           : in     vl_logic;
        ASFWRI          : in     vl_logic;
        ASFRDI          : in     vl_logic;
        OSCCLK          : in     vl_logic
    );
end ESBA;
