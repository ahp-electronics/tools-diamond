library verilog;
use verilog.vl_types.all;
entity oa_2_2 is
    port(
        A1              : in     vl_logic;
        A2              : in     vl_logic;
        B1              : in     vl_logic;
        B2              : in     vl_logic;
        Z               : out    vl_logic
    );
end oa_2_2;
