library verilog;
use verilog.vl_types.all;
entity cdr_slave_9 is
    port(
        CLK_PHASE_0     : out    vl_logic_vector(3 downto 0);
        CLK_PHASE_1     : out    vl_logic_vector(3 downto 0);
        CLK_PHASE_2     : out    vl_logic_vector(3 downto 0);
        CLK_PHASE_3     : out    vl_logic_vector(3 downto 0);
        CLK_PHASE_4     : out    vl_logic_vector(3 downto 0);
        CLK_PHASE_5     : out    vl_logic_vector(3 downto 0);
        CLK_PHASE_6     : out    vl_logic_vector(3 downto 0);
        CLK_PHASE_7     : out    vl_logic_vector(3 downto 0);
        CLK_PHASE_8     : out    vl_logic_vector(3 downto 0);
        CLKOUT_0        : out    vl_logic;
        CLKOUT_1        : out    vl_logic;
        CLKOUT_2        : out    vl_logic;
        CLKOUT_3        : out    vl_logic;
        CLKOUT_4        : out    vl_logic;
        CLKOUT_5        : out    vl_logic;
        CLKOUT_6        : out    vl_logic;
        CLKOUT_7        : out    vl_logic;
        CLKOUT_8        : out    vl_logic;
        DOUT_0          : out    vl_logic_vector(3 downto 0);
        DOUT_1          : out    vl_logic_vector(3 downto 0);
        DOUT_2          : out    vl_logic_vector(3 downto 0);
        DOUT_3          : out    vl_logic_vector(3 downto 0);
        DOUT_4          : out    vl_logic_vector(3 downto 0);
        DOUT_5          : out    vl_logic_vector(3 downto 0);
        DOUT_6          : out    vl_logic_vector(3 downto 0);
        DOUT_7          : out    vl_logic_vector(3 downto 0);
        DOUT_8          : out    vl_logic_vector(3 downto 0);
        DOUT_LOCK       : out    vl_logic_vector(8 downto 0);
        AVGING          : in     vl_logic_vector(1 downto 0);
        CLKIN_AG0_P     : in     vl_logic;
        CLKIN_AG1_P     : in     vl_logic;
        CLKIN_AG2_P     : in     vl_logic;
        CLKIN_A1_S      : in     vl_logic;
        CLKIN_A2_S      : in     vl_logic;
        CLKIN_A4_S      : in     vl_logic;
        CLKIN_A5_S      : in     vl_logic;
        CLKIN_A7_S      : in     vl_logic;
        CLKIN_A8_S      : in     vl_logic;
        CLKIN_A1_SEL    : in     vl_logic;
        CLKIN_A2_SEL    : in     vl_logic;
        CLKIN_A4_SEL    : in     vl_logic;
        CLKIN_A5_SEL    : in     vl_logic;
        CLKIN_A7_SEL    : in     vl_logic;
        CLKIN_A8_SEL    : in     vl_logic;
        CDR_LOCK_ACC    : in     vl_logic_vector(1 downto 0);
        CLK_WIDTH       : in     vl_logic;
        CDR_LOCK_MODE   : in     vl_logic;
        CIB_DATA        : in     vl_logic_vector(8 downto 0);
        CLK16           : in     vl_logic_vector(15 downto 0);
        DATA_SEL        : in     vl_logic_vector(8 downto 0);
        DIN             : in     vl_logic_vector(8 downto 0);
        EN_CLK_PHASE    : in     vl_logic;
        MASTER_LOCK     : in     vl_logic;
        OUTPUT_WIDTH    : in     vl_logic_vector(1 downto 0);
        PD_N            : in     vl_logic;
        RESET_FIFO      : in     vl_logic_vector(8 downto 0);
        RST_N           : in     vl_logic;
        TRI_ION         : in     vl_logic;
        PD_N_SLAVE      : in     vl_logic_vector(8 downto 0)
    );
end cdr_slave_9;
