library verilog;
use verilog.vl_types.all;
entity cdr_top is
    port(
        CLK_PHASE_A_0   : out    vl_logic_vector(3 downto 0);
        CLK_PHASE_A_1   : out    vl_logic_vector(3 downto 0);
        CLK_PHASE_A_2   : out    vl_logic_vector(3 downto 0);
        CLK_PHASE_D_0   : out    vl_logic_vector(3 downto 0);
        CLK_PHASE_D_1   : out    vl_logic_vector(3 downto 0);
        CLK_PHASE_D_2   : out    vl_logic_vector(3 downto 0);
        CLK_PHASE_C_0   : out    vl_logic_vector(3 downto 0);
        CLK_PHASE_C_1   : out    vl_logic_vector(3 downto 0);
        CLK_PHASE_C_2   : out    vl_logic_vector(3 downto 0);
        CLK_PHASE_B_0   : out    vl_logic_vector(3 downto 0);
        CLK_PHASE_B_1   : out    vl_logic_vector(3 downto 0);
        CLK_PHASE_B_2   : out    vl_logic_vector(3 downto 0);
        CLK_PHASE_E_0   : out    vl_logic_vector(3 downto 0);
        CLK_PHASE_E_1   : out    vl_logic_vector(3 downto 0);
        CLK_PHASE_E_2   : out    vl_logic_vector(3 downto 0);
        CLK_PHASE_F_0   : out    vl_logic_vector(3 downto 0);
        CLK_PHASE_F_1   : out    vl_logic_vector(3 downto 0);
        CLK_PHASE_F_2   : out    vl_logic_vector(3 downto 0);
        CLKOUT_A0       : out    vl_logic;
        CLKOUT_A1       : out    vl_logic;
        CLKOUT_A2       : out    vl_logic;
        CLKOUT_D0       : out    vl_logic;
        CLKOUT_D1       : out    vl_logic;
        CLKOUT_D2       : out    vl_logic;
        CLKOUT_C0       : out    vl_logic;
        CLKOUT_C1       : out    vl_logic;
        CLKOUT_C2       : out    vl_logic;
        CLKOUT_B0       : out    vl_logic;
        CLKOUT_B1       : out    vl_logic;
        CLKOUT_B2       : out    vl_logic;
        CLKOUT_E0       : out    vl_logic;
        CLKOUT_E1       : out    vl_logic;
        CLKOUT_E2       : out    vl_logic;
        CLKOUT_F0       : out    vl_logic;
        CLKOUT_F1       : out    vl_logic;
        CLKOUT_F2       : out    vl_logic;
        DOUT_A0         : out    vl_logic_vector(3 downto 0);
        DOUT_A1         : out    vl_logic_vector(3 downto 0);
        DOUT_A2         : out    vl_logic_vector(3 downto 0);
        DOUT_D0         : out    vl_logic_vector(3 downto 0);
        DOUT_D1         : out    vl_logic_vector(3 downto 0);
        DOUT_D2         : out    vl_logic_vector(3 downto 0);
        DOUT_C0         : out    vl_logic_vector(3 downto 0);
        DOUT_C1         : out    vl_logic_vector(3 downto 0);
        DOUT_C2         : out    vl_logic_vector(3 downto 0);
        DOUT_B0         : out    vl_logic_vector(3 downto 0);
        DOUT_B1         : out    vl_logic_vector(3 downto 0);
        DOUT_B2         : out    vl_logic_vector(3 downto 0);
        DOUT_E0         : out    vl_logic_vector(3 downto 0);
        DOUT_E1         : out    vl_logic_vector(3 downto 0);
        DOUT_E2         : out    vl_logic_vector(3 downto 0);
        DOUT_F0         : out    vl_logic_vector(3 downto 0);
        DOUT_F1         : out    vl_logic_vector(3 downto 0);
        DOUT_F2         : out    vl_logic_vector(3 downto 0);
        LOCKED_A0       : out    vl_logic;
        LOCKED_A1       : out    vl_logic;
        LOCKED_A2       : out    vl_logic;
        LOCKED_D0       : out    vl_logic;
        LOCKED_D1       : out    vl_logic;
        LOCKED_D2       : out    vl_logic;
        LOCKED_C0       : out    vl_logic;
        LOCKED_C1       : out    vl_logic;
        LOCKED_C2       : out    vl_logic;
        LOCKED_B0       : out    vl_logic;
        LOCKED_B1       : out    vl_logic;
        LOCKED_B2       : out    vl_logic;
        LOCKED_E0       : out    vl_logic;
        LOCKED_E1       : out    vl_logic;
        LOCKED_E2       : out    vl_logic;
        LOCKED_F0       : out    vl_logic;
        LOCKED_F1       : out    vl_logic;
        LOCKED_F2       : out    vl_logic;
        MASTER_LOCK     : out    vl_logic;
        TEST_CLK        : out    vl_logic;
        DIN_A2_CIB      : in     vl_logic;
        DIN_A1_CIB      : in     vl_logic;
        DIN_A0_CIB      : in     vl_logic;
        DIN_B2_CIB      : in     vl_logic;
        DIN_B1_CIB      : in     vl_logic;
        DIN_B0_CIB      : in     vl_logic;
        DIN_C2_CIB      : in     vl_logic;
        DIN_C1_CIB      : in     vl_logic;
        DIN_C0_CIB      : in     vl_logic;
        DIN_D2_CIB      : in     vl_logic;
        DIN_D1_CIB      : in     vl_logic;
        DIN_D0_CIB      : in     vl_logic;
        DIN_E2_CIB      : in     vl_logic;
        DIN_E1_CIB      : in     vl_logic;
        DIN_E0_CIB      : in     vl_logic;
        DIN_F2_CIB      : in     vl_logic;
        DIN_F1_CIB      : in     vl_logic;
        DIN_F0_CIB      : in     vl_logic;
        CLKIN_A_P       : in     vl_logic;
        CLKIN_D_P       : in     vl_logic;
        CLKIN_C_P       : in     vl_logic;
        CLKIN_A1_S      : in     vl_logic;
        CLKIN_A2_S      : in     vl_logic;
        CLKIN_D1_S      : in     vl_logic;
        CLKIN_D2_S      : in     vl_logic;
        CLKIN_C1_S      : in     vl_logic;
        CLKIN_C2_S      : in     vl_logic;
        CLKIN_B_P       : in     vl_logic;
        CLKIN_E_P       : in     vl_logic;
        CLKIN_F_P       : in     vl_logic;
        CLKIN_B1_S      : in     vl_logic;
        CLKIN_B2_S      : in     vl_logic;
        CLKIN_E1_S      : in     vl_logic;
        CLKIN_E2_S      : in     vl_logic;
        CLKIN_F1_S      : in     vl_logic;
        CLKIN_F2_S      : in     vl_logic;
        DIN_A0_PAD      : in     vl_logic;
        DIN_A1_PAD      : in     vl_logic;
        DIN_A2_PAD      : in     vl_logic;
        DIN_D0_PAD      : in     vl_logic;
        DIN_D1_PAD      : in     vl_logic;
        DIN_D2_PAD      : in     vl_logic;
        DIN_C0_PAD      : in     vl_logic;
        DIN_C1_PAD      : in     vl_logic;
        DIN_C2_PAD      : in     vl_logic;
        DIN_B0_PAD      : in     vl_logic;
        DIN_B1_PAD      : in     vl_logic;
        DIN_B2_PAD      : in     vl_logic;
        DIN_E0_PAD      : in     vl_logic;
        DIN_E1_PAD      : in     vl_logic;
        DIN_E2_PAD      : in     vl_logic;
        DIN_F0_PAD      : in     vl_logic;
        DIN_F1_PAD      : in     vl_logic;
        DIN_F2_PAD      : in     vl_logic;
        MC1_EN_TEST_CLK : in     vl_logic;
        MC1_EN_CLK_PHASE_ADC: in     vl_logic;
        MC1_EN_CLK_PHASE_BEF: in     vl_logic;
        MC1_ALU_BW      : in     vl_logic_vector(1 downto 0);
        MC1_AVGING_ADC  : in     vl_logic_vector(1 downto 0);
        MC1_AVGING_BEF  : in     vl_logic_vector(1 downto 0);
        MC1_CDR_LOCKACC_ADC: in     vl_logic_vector(1 downto 0);
        MC1_CDR_LOCKACC_BEF: in     vl_logic_vector(1 downto 0);
        MC1_CDR_LOCKMODE_ADC: in     vl_logic;
        MC1_CDR_LOCKMODE_BEF: in     vl_logic;
        MC1_DOUT_CLKIN_SEL_A1: in     vl_logic;
        MC1_DOUT_CLKIN_SEL_B1: in     vl_logic;
        MC1_DOUT_CLKIN_SEL_A2: in     vl_logic;
        MC1_DOUT_CLKIN_SEL_B2: in     vl_logic;
        MC1_DOUT_CLKIN_SEL_D1: in     vl_logic;
        MC1_DOUT_CLKIN_SEL_E1: in     vl_logic;
        MC1_DOUT_CLKIN_SEL_D2: in     vl_logic;
        MC1_DOUT_CLKIN_SEL_E2: in     vl_logic;
        MC1_DOUT_CLKIN_SEL_C1: in     vl_logic;
        MC1_DOUT_CLKIN_SEL_F1: in     vl_logic;
        MC1_DOUT_CLKIN_SEL_C2: in     vl_logic;
        MC1_DOUT_CLKIN_SEL_F2: in     vl_logic;
        MC1_REFCLK_SEL  : in     vl_logic;
        MC1_DIN_SEL_A0  : in     vl_logic;
        MC1_DIN_SEL_A1  : in     vl_logic;
        MC1_DIN_SEL_A2  : in     vl_logic;
        MC1_DIN_SEL_B0  : in     vl_logic;
        MC1_DIN_SEL_B1  : in     vl_logic;
        MC1_DIN_SEL_B2  : in     vl_logic;
        MC1_DIN_SEL_C0  : in     vl_logic;
        MC1_DIN_SEL_C1  : in     vl_logic;
        MC1_DIN_SEL_C2  : in     vl_logic;
        MC1_DIN_SEL_D0  : in     vl_logic;
        MC1_DIN_SEL_D1  : in     vl_logic;
        MC1_DIN_SEL_D2  : in     vl_logic;
        MC1_DIN_SEL_E0  : in     vl_logic;
        MC1_DIN_SEL_E1  : in     vl_logic;
        MC1_DIN_SEL_E2  : in     vl_logic;
        MC1_DIN_SEL_F0  : in     vl_logic;
        MC1_DIN_SEL_F1  : in     vl_logic;
        MC1_DIN_SEL_F2  : in     vl_logic;
        FORCE_LOCK      : in     vl_logic;
        MASTER_HOLD     : in     vl_logic;
        MC1_OUTPUT_WIDTH_ADC: in     vl_logic_vector(1 downto 0);
        MC1_OUTPUT_WIDTH_BEF: in     vl_logic_vector(1 downto 0);
        MC1_PD_N_ADC    : in     vl_logic;
        MC1_PD_N_BEF    : in     vl_logic;
        MC1_PD_N        : in     vl_logic;
        MC1_REFLOCK_ACC : in     vl_logic_vector(1 downto 0);
        MC1_FIFO_BYPASS_A: in     vl_logic_vector(2 downto 0);
        MC1_FIFO_BYPASS_D: in     vl_logic_vector(2 downto 0);
        MC1_FIFO_BYPASS_C: in     vl_logic_vector(2 downto 0);
        MC1_FIFO_BYPASS_B: in     vl_logic_vector(2 downto 0);
        MC1_FIFO_BYPASS_E: in     vl_logic_vector(2 downto 0);
        MC1_FIFO_BYPASS_F: in     vl_logic_vector(2 downto 0);
        MC1_SEL_WIDTH   : in     vl_logic;
        MC1_TEST_CLK_SEL: in     vl_logic_vector(3 downto 0);
        REFCLK_EDGE     : in     vl_logic;
        REFCLK_PRIM     : in     vl_logic;
        MACO_RST_N      : in     vl_logic;
        TRI_ION         : in     vl_logic;
        RSTN            : in     vl_logic;
        RSTN_A2         : in     vl_logic;
        RSTN_A1         : in     vl_logic;
        RSTN_A0         : in     vl_logic;
        RSTN_B2         : in     vl_logic;
        RSTN_B1         : in     vl_logic;
        RSTN_B0         : in     vl_logic;
        RSTN_C2         : in     vl_logic;
        RSTN_C1         : in     vl_logic;
        RSTN_C0         : in     vl_logic;
        RSTN_D2         : in     vl_logic;
        RSTN_D1         : in     vl_logic;
        RSTN_D0         : in     vl_logic;
        RSTN_E2         : in     vl_logic;
        RSTN_E1         : in     vl_logic;
        RSTN_E0         : in     vl_logic;
        RSTN_F2         : in     vl_logic;
        RSTN_F1         : in     vl_logic;
        RSTN_F0         : in     vl_logic;
        MC1_GSRN_EN     : in     vl_logic
    );
end cdr_top;
