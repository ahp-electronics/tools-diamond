library verilog;
use verilog.vl_types.all;
entity flash_qual is
    port(
        fl_init_addr_cfg_exec_a: out    vl_logic;
        fl_init_addr_trim_exec_a: out    vl_logic;
        fl_init_addr_fea_exec_a: out    vl_logic;
        fl_init_addr_ufm_exec_a: out    vl_logic;
        fl_write_addr_exec_a: out    vl_logic;
        fl_prog_incr_nv_exec_a: out    vl_logic;
        fl_prog_tag_exec_a: out    vl_logic;
        fl_prog_udss_exec_a: out    vl_logic;
        fl_prog_ufs_exec_a: out    vl_logic;
        fl_prog_trim_exec_a: out    vl_logic_vector(5 downto 0);
        fl_prog_feat_exec_a: out    vl_logic_vector(5 downto 0);
        fl_read_incr_nv_exec_a: out    vl_logic;
        fl_read_tag_exec_a: out    vl_logic;
        fl_read_trim3_exec_a: out    vl_logic;
        fl_mtest_exec_a : out    vl_logic;
        sector_dat_a    : out    vl_logic_vector(7 downto 0);
        exec_buf_reset_a: out    vl_logic;
        fl_prog_64_exec_a: out    vl_logic;
        fl_exec_buf_a   : in     vl_logic_vector(127 downto 0);
        exec_buf_ready_a: in     vl_logic;
        sect_cfg_sel_a  : in     vl_logic;
        sect_ufm_sel_a  : in     vl_logic;
        sect_trim_sel_a : in     vl_logic;
        sect_feat_sel_a : in     vl_logic;
        sec_row_active_a: in     vl_logic;
        trim_row4_active_a: in     vl_logic;
        fl_init_addr_cfg_exec_b: out    vl_logic;
        fl_init_addr_trim_exec_b: out    vl_logic;
        fl_init_addr_fea_exec_b: out    vl_logic;
        fl_init_addr_ufm_exec_b: out    vl_logic;
        fl_write_addr_exec_b: out    vl_logic;
        fl_prog_incr_nv_exec_b: out    vl_logic;
        fl_prog_tag_exec_b: out    vl_logic;
        fl_prog_udss_exec_b: out    vl_logic;
        fl_prog_ufs_exec_b: out    vl_logic;
        fl_prog_trim_exec_b: out    vl_logic_vector(5 downto 0);
        fl_prog_feat_exec_b: out    vl_logic_vector(5 downto 0);
        fl_read_incr_nv_exec_b: out    vl_logic;
        fl_read_tag_exec_b: out    vl_logic;
        fl_read_trim3_exec_b: out    vl_logic;
        fl_mtest_exec_b : out    vl_logic;
        sector_dat_b    : out    vl_logic_vector(7 downto 0);
        exec_buf_reset_b: out    vl_logic;
        fl_prog_64_exec_b: out    vl_logic;
        fl_exec_buf_b   : in     vl_logic_vector(127 downto 0);
        exec_buf_ready_b: in     vl_logic;
        sect_cfg_sel_b  : in     vl_logic;
        sect_ufm_sel_b  : in     vl_logic;
        sect_trim_sel_b : in     vl_logic;
        sect_feat_sel_b : in     vl_logic;
        sec_row_active_b: in     vl_logic;
        trim_row4_active_b: in     vl_logic;
        fl_init_addr_cfg_exec_c: out    vl_logic;
        fl_init_addr_trim_exec_c: out    vl_logic;
        fl_init_addr_fea_exec_c: out    vl_logic;
        fl_init_addr_ufm_exec_c: out    vl_logic;
        fl_write_addr_exec_c: out    vl_logic;
        fl_prog_incr_nv_exec_c: out    vl_logic;
        fl_prog_tag_exec_c: out    vl_logic;
        fl_prog_udss_exec_c: out    vl_logic;
        fl_prog_ufs_exec_c: out    vl_logic;
        fl_prog_trim_exec_c: out    vl_logic_vector(5 downto 0);
        fl_prog_feat_exec_c: out    vl_logic_vector(5 downto 0);
        fl_read_incr_nv_exec_c: out    vl_logic;
        fl_read_tag_exec_c: out    vl_logic;
        fl_read_trim3_exec_c: out    vl_logic;
        fl_mtest_exec_c : out    vl_logic;
        sector_dat_c    : out    vl_logic_vector(7 downto 0);
        exec_buf_reset_c: out    vl_logic;
        fl_prog_64_exec_c: out    vl_logic;
        fl_exec_buf_c   : in     vl_logic_vector(127 downto 0);
        exec_buf_ready_c: in     vl_logic;
        sect_cfg_sel_c  : in     vl_logic;
        sect_ufm_sel_c  : in     vl_logic;
        sect_trim_sel_c : in     vl_logic;
        sect_feat_sel_c : in     vl_logic;
        sec_row_active_c: in     vl_logic;
        trim_row4_active_c: in     vl_logic;
        isc_rst_async   : in     vl_logic;
        isc_rst_sync    : in     vl_logic;
        smclk           : in     vl_logic;
        mfg_flash_en    : in     vl_logic;
        access_sudo     : in     vl_logic;
        fl_erase_qual   : in     vl_logic;
        fl_erase_all_qual: in     vl_logic;
        fl_prog_ucode_qual: in     vl_logic;
        fl_prog_done_qual: in     vl_logic;
        fl_prog_sec_qual: in     vl_logic;
        fl_prog_secplus_qual: in     vl_logic;
        fl_disable_done0_qual: in     vl_logic;
        fl_disable_done1_qual: in     vl_logic;
        fl_prog_authmode_qual: in     vl_logic;
        fl_prog_aesfea_qual: in     vl_logic;
        fl_init_addr_qual: in     vl_logic;
        fl_write_addr_qual: in     vl_logic;
        fl_prog_incr_nv_qual: in     vl_logic;
        fl_read_incr_nv_qual: in     vl_logic;
        fl_prog_password_qual: in     vl_logic;
        fl_prog_feature_qual: in     vl_logic;
        fl_prog_feabits_qual: in     vl_logic;
        fl_init_addr_ufm_qual: in     vl_logic;
        fl_prog_tag_qual: in     vl_logic;
        fl_erase_tag_qual: in     vl_logic;
        fl_read_tag_qual: in     vl_logic;
        fl_prog_pes_qual: in     vl_logic;
        fl_prog_mes_qual: in     vl_logic;
        fl_prog_hes_qual: in     vl_logic;
        fl_prog_trim0_qual: in     vl_logic;
        fl_prog_trim1_qual: in     vl_logic;
        fl_read_hes_qual: in     vl_logic;
        fl_mtest_qual   : in     vl_logic;
        fl_prog_pubkey0_qual: in     vl_logic;
        fl_prog_pubkey1_qual: in     vl_logic;
        fl_prog_pubkey2_qual: in     vl_logic;
        fl_prog_pubkey3_qual: in     vl_logic;
        fl_prog_aeskey0_qual: in     vl_logic;
        fl_prog_aeskey1_qual: in     vl_logic;
        fl_prog_usec_qual: in     vl_logic;
        fl_prog_csec_qual: in     vl_logic;
        fl_prog_uds_qual: in     vl_logic;
        fl_busy_all     : in     vl_logic;
        fl_exec_buf     : out    vl_logic_vector(127 downto 0);
        current_sector  : out    vl_logic_vector(11 downto 0);
        sector_dat      : in     vl_logic_vector(15 downto 0);
        isc_exec_e      : in     vl_logic;
        blk_sel         : in     vl_logic_vector(1 downto 0);
        sector_erase    : in     vl_logic_vector(11 downto 0);
        mfg_fl_pp       : in     vl_logic;
        mfg_mtest_fl_sel: in     vl_logic_vector(1 downto 0)
    );
end flash_qual;
