--
@ER--B$FbsEHo0OR52gR4g-cRRj.jd$R1MHbDO$H0ROQM
R--fN]C8:CsR#//$DMbH0OH$N/lb..jjDjdNl0/NCbbsG#/HMDHGH/DLC/oMHCsOC/oMC_oMHCsOs./N_lMsPI3E48yR-f
--

--
-
R--1bHlD)CRqIvRHR0E#oHMDqCR7 7)1V1RFLsRFR0Es8CNR8NMRHIs0-C
-NRas0oCRX:RHMDHGD

HNLssH$RC;CC
#
kCCRHC#C30D8_FOoH_n44cD3NDk;
#HCRC3CC#_08DHFoOH_#o8MC3DND;H
DLssN$MRkHl#H;#
kCMRkHl#H3FPOlMbFC#M03DND;M
C0$H0Rv)qhW_)R
H#RRRRoCCMsRHO5R
RRRRRRNRVl$HDR#:R0MsHo=R:RF"MM;C"
RRRRRRRR8IH0:ERR0HMCsoCRR:=4Rj;
RRRRRRRR8N8s8IH0:ERR0HMCsoCRR:=4Rd;RRRRR-RR-HRLoMRCFEkoRsVFRb8C0RE
RRRRR8RRCEb0RH:RMo0CC:sR=4RUg
.;RRRRRRRR80Fk_osCRL:RFCFDN:MR=NRVD;#CRRRRRR--ERN#Fbk0ks0RCRo
RRRRR8RRHsM_C:oRRFLFDMCNRR:=V#NDCR;RRRRR-E-RN8#RNR0NHkMb0CRsoR
SRsRR#80_NR0N:0R#soHM;S
SIls_FR8C:0R#soHMRR:="QW)aw _Qa)1"R;
RRRRRNRR8_8ssRCo:FRLFNDCM=R:Rk0sCRRRR-RR-NRE88RN8#sC#CRsoR
RRRRRR;R2
RRRRsbF0
R5RRRRRRRR7amz:kRF00R#8F_Do_HOP0COFIs5HE80-84RF0IMF2Rj;R
RRRRRRQR7h:RRRRHM#_08DHFoOC_POs0F58IH04E-RI8FMR0Fj
2;RRRRRRRRq)77RH:RM0R#8F_Do_HOP0COFNs58I8sHE80-84RF0IMF2Rj;R
RRRRRR RWRRR:H#MR0D8_FOoH;RRRRRRR-I-RsCH0RNCMLRDCVRFss
NlRRRRRRRRBRpi:MRHR8#0_oDFHRO;RRRRR-R-RFODOV	RFssRNRl,Ns88,HR8MS
SmiBpRH:RM0R#8F_Do;HO
)SS1:aRRRHM#_08DHFoOR;RRRRRRR--sCC#0MRFR0FkbRk0s
CoShS RH:RM0R#8F_DoSHOS-RR-MRCRMbHRRFVLODF	NRslS
S2C;
MC8RM00H$qR)v)h_W
;
NEsOHO0C0CksRFLDOs	_NFlRVqR)v)h_W#RH
MVkOF0HMkRVMHO_M5H0LRR:LDFFC2NMR0sCkRsM#H0sMHoR#C
Lo
HMRVRHR25LRC0EMR
RRCRs0Mks52"";R
RCCD#
RRRR0sCk5sM"kBFDM8RFH0RlCbDl0CMRFADO)	RqRv3Q0#REsCRCRN8Ns88CR##sHCo#s0CCk8R#oHMRC0ERl#NCDROFRO	N0#RE)CRq"v?2R;
R8CMR;HV
8CMRMVkOM_HH
0;Ns00H0LkCCRoMNCs0_FssFCbs:0RRs#0H;Mo
N--0H0sLCk0RMoCC0sNFss_CsbF0VRFRFLDOs	_N:lRRONsECH0Os0kC#RHRMVkOM_HH805F_k0s2Co;k
VMHO0F#MR0MsHoD.#PR5N:0R#soHM2CRs0MksR8#0_oDFHPO_CFO0s#RH
sPNHDNLCDR#PRR:#_08DHFoOC_POs0F5EN'H-oENF'DIFR8IFM0R;j2
sPNHDNLCRRH:MRH0CCosL;
CMoH
VRRFHsRRRHMjFR0RP#D'oEHEFRDFRb
RHRRVNR55EN'H-oEH=2RR''42ER0CSM
RDR#P25HRR:=';4'
DSC#SC
RDR#P25HRR:=';j'
MSC8VRH;R
RCRM8DbFF;R
RskC0s#MRD
P;CRM8#H0sM#o.D
P;VOkM0MHFRP#D.s#0H5MoNRR:#_08DHFoOC_POs0F2CRs0MksRs#0HRMoHP#
NNsHLRDC#RR:#H0sMNo5'oEHE'-ND+FI4FR8IFM0R;42
sPNHDNLCRRH:MRH0CCosL;
CMoH
VRRFHsRRRHMNF'DIFR0REN'HRoEDbFF
RRRRRHV5HN52RR='24'RC0EMR
SRH#5-DN'F4I+2=R:R''4;C
SD
#CS#RR5NH-'IDF+R42:'=Rj
';S8CMR;HV
CRRMD8RF;Fb
sRRCs0kM;R#
8CMRP#D.s#0H;Mo
0N0skHL0GCROs_bFRb#:0R#soHM;-
-O#FM00NMRP#sN:DRR8#0_oDFHPO_CFO0sH5I8-0E4FR8IFM0RRj2:#=R0MsHoD.#P#5s0N_80;N2
R--LHCoMDRLFRO	sRNlHDlbCMlC0HN0F#MRHNoMDV#
k0MOHRFMo_C0OHEFOIC_HE8058IH0:ERR0HMCsoC2CRs0MksR0HMCsoCR
H#PHNsNCLDRDPNRH:RMo0CC:sR=;Rj
sPNHDNLCHR8P,d.RP8H4Rn,8UHP,HR8PRc,8.HP,HR8P:4RR0HMCsoC;C
Lo
HMRHR8PRd.:5=RI0H8E2-4/;dn
8RRHnP4RR:=58IH04E-2U/4;R
R8UHPRR:=58IH04E-2;/g
8RRHRPc:5=RI0H8E2-4/
c;RHR8P:.R=IR5HE80-/42.R;
RP8H4=R:RH5I8-0E4
2;RVRHRH58P>4RRRj20MEC
RRRRDPNRR:=PRND+;R4
CRRMH8RVR;
RRHV5P8H.RR>j02RE
CMRRRRPRND:P=RN+DRR
4;RMRC8VRH;R
RH5VR8cHPRj>R2ER0CRM
RPRRN:DR=NRPDRR+4R;
R8CMR;HV
HRRV8R5HRPU>2RjRC0EMR
RRNRPD=R:RDPNR4+R;R
RCRM8H
V;RVRHRH58PR4n>2RjRC0EMR
RRNRPD=R:RDPNR4+R;R
RCRM8H
V;-R-RH5VR8dHP.RR>j02RE
CM-R-RRNRPD=R:RDPNR4+R;-
-RMRC8VRH;R
RH5VRPRND>2R.RC0EMR
RRCRs0MksRR5.*P*RN+DRR*.R*PR5N-DRR2d2;R
RCCD#
RRRR0sCkRsM5*.R*NRPD
2;RMRC8VRH;RRRRRRR
8CMR0oC_FOEH_OCI0H8EV;
k0MOHRFMo_C0OHEFO8C_CEb05b8C0:ERR0HMCsoC2CRs0MksR0HMCsoCR
H#PHNsNCLDRO8_EOFHCC_8bR0E:MRH0CCos=R:R
j;LHCoMR
RH5VR80CbERR>U.4g2ER0CRM
R8RR_FOEH_OC80CbE=R:Rd4nU
c;RDRC#RHV5b8C0<ER=4RUgN.RM88RCEb0Rc>RjRgn2ER0CRM
R8RR_FOEH_OC80CbE=R:RgU4.R;
R#CDH5VR80CbE=R<RgcjnMRN8CR8bR0E>jR.cRU20MEC
RRRRO8_EOFHCC_8bR0E:c=Rj;gn
CRRDV#HRC58bR0E<.=RjRcUNRM880CbERR>4cj.R02RE
CMRRRR8E_OFCHO_b8C0:ER=jR.c
U;RDRC#RHV5b8C0<ER=jR4.NcRM88RCEb0R6>R4R.20MEC
RRRRO8_EOFHCC_8bR0E:4=Rj;.c
CRRDV#HRC58bR0E<6=R4R.20MEC
RRRRO8_EOFHCC_8bR0E:6=R4
.;RMRC8VRH;R
RskC0s8MR_FOEH_OC80CbEC;
Mo8RCO0_EOFHCC_8b;0E
MVkOF0HMCRo0H_I8_0El_F8UE5OFCHO_RI8:MRH0CCoss2RCs0kMMRH0CCos#RH
sPNHDNLCHRI8_0El_F8URR:HCM0o;Cs
oLCHRM
RRHV5FOEH_OCI>8RRRU20MEC
RRRR8IH0lE_FU8_RR:=OHEFOIC_8RR-5FOEH_OCIl8RFU8R2R;
R#CDCR
RRHRI8_0El_F8U=R:RFOEH_OCI
8;RMRC8VRH;R
RskC0sIMRHE80_8lF_
U;CRM8o_C0I0H8EF_l8;_U
F
OMN#0MI0R_FOEH_OCI0H8ERR:HCM0oRCs:o=RCO0_EOFHCH_I850EI0H8E
2;O#FM00NMROI_EOFHCC_8bR0E:MRH0CCos=R:Rd4nUoc/CI0_HE80_8lF_IU5_FOEH_OCI0H8E
2;O#FM00NMRO8_EOFHCC_8bR0E:MRH0CCos=R:R0oC_FOEH_OC80CbEC58b20E;F
OMN#0M80R_FOEH_OCI0H8ERR:HCM0oRCs:5=R4Undc_/8OHEFO8C_CEb02RR+5n54d/Uc8E_OFCHO_b8C0RE2/2RU;V

k0MOHRFMo_C0M_klODCD#85IRH:RMo0CCOs;EOFHC8_IRH:RMo0CCRs2skC0sHMRMo0CCHsR#N
PsLHNDMCRkOl_C#DDRH:RMo0CC
s;LHCoMR
RM_klODCD#=R:R85I-/42OHEFOIC_8RR+4R;
R0sCkRsMM_klODCD#C;
Mo8RCM0_kOl_C#DD;V

k0MOHRFMo_C0#CHx5OIMRH:RMo0CCRs;8RMO:MRH0CCoss2RCs0kMMRH0CCos#RH
oLCHRM
RCRs0MksROIMR8*RM
O;CRM8o_C0#CHx;V

k0MOHRFMo_C0LDFF8_58#CHxRH:RMo0CCRs;IH_#x:CRR0HMCsoC;_R8O:IRR0HMCsoC;_RIO:IRR0HMCsoC2CRs0MksR0HMCsoCR
H#LHCoMV
HR_58#CHxRR<=IH_#xRC20MEC
sRRCs0kM_R8O
I;CCD#
sRRCs0kM_RIO
I;CRM8H
V;CRM8o_C0LDFF8V;
k0MOHRFMo_C0C_M880CbEH5#x:CRR0HMCsoCR8;RCEb0RH:RMo0CCRs2skC0sHMRMo0CCHsR#N
PsLHNDlCRH#M_HRxC:MRH0CCos=R:R
j;LHCoMR
Rl_HM#CHxRR:=80CbER;
RRHV5x#HCRR<80CbE02RE
CMRRRRl_HM#CHxRR:=#CHx;R
RCRM8H
V;RCRs0MksRMlH_x#HCC;
Mo8RCC0_M88_CEb0;O

F0M#NRM0OHEFOIC_HE80RH:RMo0CC:sR=CRo0F_LF5D8o_C0#CHx50oC_lMk_DOCDI#5HE80,_R8OHEFOIC_HE802C,o0k_MlC_OD5D#80CbE8,R_FOEH_OC80CbE,22
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRCRo0H_#xoC5CM0_kOl_C#DD58IH0RE,IE_OFCHO_8IH0,E2o_C0M_klODCD#C58b,0EROI_EOFHCC_8b20E2S,
SSSSSSSSS8SR_FOEH_OCI0H8EI,R_FOEH_OCI0H8E
2;O#FM00NMR8IH0ME_kOl_C#DDRH:RMo0CC:sR=CRo0F_LF5D8o_C0#CHx50oC_lMk_DOCDI#5HE80,_R8OHEFOIC_HE802C,o0k_MlC_OD5D#80CbE8,R_FOEH_OC80CbE,22
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR0oC_x#HCC5o0k_MlC_OD5D#I0H8EI,R_FOEH_OCI0H8Eo2,CM0_kOl_C#DD5b8C0RE,IE_OFCHO_b8C02E2,S
SSSSSSSSSSRRRRH5I8-0E482/_FOEH_OCI0H8E5,RI0H8E2-4/OI_EOFHCH_I820ER4+R;F
OMN#0M80RCEb0_lMk_DOCD:#RR0HMCsoCRR:=o_C0LDFF8C5o0H_#xoC5CM0_kOl_C#DD58IH0RE,8E_OFCHO_8IH0,E2o_C0M_klODCD#C58b,0ERO8_EOFHCC_8b20E2R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRCRo0H_#xoC5CM0_kOl_C#DD58IH0RE,IE_OFCHO_8IH0,E2o_C0M_klODCD#C58b,0EROI_EOFHCC_8b20E2S,
SSSSSSSSSRRR5b8C04E-2_/8OHEFO8C_CEb0,8R5CEb0-/42IE_OFCHO_b8C0RE2+;R4SOR
F0M#NRM0xFCsR#:R0D8_FOoH_OPC05FsOHEFOIC_HE80*8IH0ME_kOl_C#DD-8IH04E-RI8FMR0Fj:2R=FR50sEC#>R=R''j2O;
F0M#NRM0#NsPDD_#PRR:#_08DHFoOC_POs0F5FOEH_OCI0H8EH*I8_0EM_klODCD#R-48MFI0jFR2=R:RsxCFRR&#H0sM#o.DsP5#80_N20N;F
OMN#0M#0RsDPNR#:R0MsHoE5OFCHO_8IH0IE*HE80_lMk_DOCD8#RF0IMF2R4RR:=#.DP#H0sM#o5sDPN_P#D2-;
-o#HM#NDRsVFRMMF-ED#N8bCRFLDOs	RN
l#0C$bR0Fk_#Lk4$_0bHCR#sRNsRN$5b8C0ME_kOl_C#DD-84RF0IMF,RjR8IH0ME_kOl_C#DD-84RF0IMF2RjRRFV#_08DHFoO#;
HNoMDkRF0k_L#:4RR0Fk_#Lk4$_0bRC;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-7R.RsNsNF$RVFR8k50RHkMb0FR0RH0s-N#002C#
b0$CkRF0k_L#0._$RbCHN#Rs$sNRC58b_0EM_klODCD#R-48MFI0jFR,*R.I0H8Ek_MlC_OD+D#4FR8IFM0RRj2F#VR0D8_FOoH;H
#oDMNR0Fk_#Lk.RR:F_k0L.k#_b0$CR;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RR.7NNss$VRFRk8F0HR5M0bkRR0F0-sH#00NC
#20C$bR0Fk_#Lkc$_0bHCR#sRNsRN$5b8C0ME_kOl_C#DD-84RF0IMF,RjRIc*HE80_lMk_DOCDd#+RI8FMR0FjF2RV0R#8F_Do;HO
o#HMRNDF_k0Lck#RF:RkL0_k_#c0C$b;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--.N7Rs$sNRRFV80FkRM5HbRk000FRs#H-0CN0#02
$RbCF_k0LUk#_b0$C#RHRsNsN5$R80CbEk_MlC_OD-D#4FR8IFM0RRj,UH*I8_0EM_klODCD#R+(8MFI0jFR2VRFR8#0_oDFH
O;#MHoNFDRkL0_kR#U:kRF0k_L#0U_$;bCRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-.-R7sRNsRN$F8VRFRk05bHMk00RFsR0H0-#N#0C2$
0bbCRN0sH$k_L#0U_$RbCHN#Rs$sNRC58b_0EM_klODCD#R-48MFI0jFR,HRI8_0EM_klODCD#R-48MFI0jFR2VRFR8#0_oDFH
O;#MHoNbDRN0sH$k_L#:URRsbNH_0$LUk#_b0$CR;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-.-R7sRNsRN$F8VRFRk05bHMk00RFsR0H0-#N#0C2$
0bFCRkL0_kn#4_b0$C#RHRsNsN5$R80CbEk_MlC_OD-D#4FR8IFM0RRj,4In*HE80_lMk_DOCD4#+6FR8IFM0RRj2F#VR0D8_FOoH;H
#oDMNR0Fk_#Lk4:nRR0Fk_#Lk40n_$;bCRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RR.7NNss$VRFRk8F0HR5M0bkRR0F0-sH#00NC
#20C$bRsbNH_0$L4k#n$_0bHCR#sRNsRN$5b8C0ME_kOl_C#DD-84RF0IMF,RjRI.*HE80_lMk_DOCD4#+RI8FMR0FjF2RV0R#8F_Do;HO
o#HMRNDbHNs0L$_kn#4Rb:RN0sH$k_L#_4n0C$b;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--.N7Rs$sNRRFV80FkRM5HbRk000FRs#H-0CN0#02
$RbCF_k0Ldk#.$_0bHCR#sRNsRN$5b8C0ME_kOl_C#DD-84RF0IMF,RjR*d.I0H8Ek_MlC_OD+D#d84RF0IMF2RjRRFV#_08DHFoO#;
HNoMDkRF0k_L#Rd.:kRF0k_L#_d.0C$b;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-7R.RsNsNF$RVFR8k50RHkMb0FR0RH0s-N#002C#
b0$CNRbs$H0_#Lkd0._$RbCHN#Rs$sNRC58b_0EM_klODCD#R-48MFI0jFR,*RcI0H8Ek_MlC_OD+D#dFR8IFM0RRj2F#VR0D8_FOoH;H
#oDMNRsbNH_0$Ldk#.RR:bHNs0L$_k.#d_b0$CR;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RR.7NNss$VRFRk8F0HR5M0bkRR0F0-sH#00NC
#2#MHoNFDRkC0_MRR:#_08DHFoOC_POs0F5b8C0ME_kOl_C#DD-84RF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RNCML#DCRsVFRH0s-N#00
C##MHoNIDRsC0_MRR:#_08DHFoOC_POs0F5b8C0ME_kOl_C#DD-84RF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RHIs0CCRMDNLCV#RFCsRNROEsRFIF)VRqOvRC#DD
o#HMRNDHsM_C:oRR8#0_oDFHPO_CFO0sH5I8+0Ed86RF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-k-R#RC80sFRC#oH0RCs7RQh
o#HMRNDF_k0sRCo:0R#8F_Do_HOP0COFIs5HE80+Rd68MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-k-R#RC80sFRC#oH0RCs7amz
o#HMRNDNs8_C:oRR8#0_oDFHPO_CFO0s85N8HsI8-0E4FR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-#RkC08RFCRso0H#CqsR7
7)#MHoNDDRFNI_8R8s:0R#8F_Do_HOP0COF4s5dFR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-8RN8LsRHR0#HkMb0FR0Rv)qRDOCD5#RcHRL0s#RCHJks2C8
o#HMRNDNC8soRR:#_08DHFoOC_POs0F58N8s8IH04E-RI8FMR0FjR2;-0-RFCRso0H#C0sRE#CRCODC0HR#oDMNRRFV0#sH0CN0
R--CRM8LODF	NRsllRHblDCCNM00MHFRo#HM#ND
0N0skHL0\CR3lsN_VFV#\C0R#:R0MsHo
;
LHCoMR
R
RRRRR--QNVR8I8sHE80RO<REOFHCH_I8R0ENH##o'MRj0'RFMRkk8#CR0LH#R
RRjRzRRR:H5VRNs88I0H8ERR=4o2RCsMCN
0CSRRRRIDF_8N8s=R<Rj"jjjjjjjjjj"jjRN&R8C_so25j;C
SMo8RCsMCNR0Cz
j;RRRRzR4R:VRHR85N8HsI8R0E=2R.RMoCC0sNCR
SRDRRFNI_8R8s<"=Rjjjjjjjjjjjj"RR&Ns8_C4o5RI8FMR0Fj
2;S8CMRMoCC0sNC4Rz;R
RR.RzRRR:H5VRNs88I0H8ERR=do2RCsMCN
0CSRRRRIDF_8N8s=R<Rj"jjjjjjjjjj&"RR_N8s5Co.FR8IFM0R;j2
MSC8CRoMNCs0zCR.R;
RzRRd:RRRRHV58N8s8IH0=ERRRc2oCCMsCN0
RSRRFRDI8_N8<sR=jR"jjjjjjjjj&"RR_N8s5CodFR8IFM0R;j2
MSC8CRoMNCs0zCRdR;
RzRRc:RRRRHV58N8s8IH0=ERRR62oCCMsCN0
RSRRFRDI8_N8<sR=jR"jjjjjjjj"RR&Ns8_Cco5RI8FMR0Fj
2;S8CMRMoCC0sNCcRz;R
RR6RzRRR:H5VRNs88I0H8ERR=no2RCsMCN
0CSRRRRIDF_8N8s=R<Rj"jjjjjjRj"&8RN_osC586RF0IMF2Rj;C
SMo8RCsMCNR0Cz
6;RRRRzRnR:VRHR85N8HsI8R0E=2R(RMoCC0sNCR
SRDRRFNI_8R8s<"=Rjjjjj"jjRN&R8C_soR5n8MFI0jFR2S;
CRM8oCCMsCN0R;zn
RRRRRz(RH:RVNR58I8sHE80RU=R2CRoMNCs0SC
RRRRD_FINs88RR<="jjjj"jjRN&R8C_soR5(8MFI0jFR2S;
CRM8oCCMsCN0R;z(
RRRRRzURH:RVNR58I8sHE80Rg=R2CRoMNCs0SC
RRRRD_FINs88RR<="jjjjRj"&8RN_osC58URF0IMF2Rj;C
SMo8RCsMCNR0Cz
U;RRRRzRgR:VRHR85N8HsI8R0E=jR42CRoMNCs0SC
RRRRD_FINs88RR<="jjjj&"RR_N8s5CogFR8IFM0R;j2
MSC8CRoMNCs0zCRgR;
RzRR4RjR:VRHR85N8HsI8R0E=4R42CRoMNCs0SC
RRRRD_FINs88RR<="jjj"RR&Ns8_C4o5jFR8IFM0R;j2
MSC8CRoMNCs0zCR4
j;RRRRzR44RH:RVNR58I8sHE80R4=R.o2RCsMCN
0CSRRRRIDF_8N8s=R<Rj"j"RR&Ns8_C4o54FR8IFM0R;j2
MSC8CRoMNCs0zCR4
4;RRRRzR4.RH:RVNR58I8sHE80R4=Rdo2RCsMCN
0CSRRRRIDF_8N8s=R<R''jRN&R8C_so.54RI8FMR0Fj
2;S8CMRMoCC0sNC4Rz.R;
RzRR4RdR:VRHR85N8HsI8R0E>dR42CRoMNCs0SC
RRRRD_FINs88RR<=Ns8_C4o5dFR8IFM0R;j2
MSC8CRoMNCs0zCR4
d;
RRRRR--Q5VR8_HMs2CoRosCHC#0sQR7h#RkHRMoB
piRRRRzR4cRH:RV8R5HsM_CRo2oCCMsCN0
RRRRRRRRFbsO#C#Rp5Bi7,RQRh2LHCoMR
RRRRRRRRRRVRHRp5BiRR='R4'NRM8B'piCMPC002RE
CMRRRRRRRRRRRRRRRRHsM_C<oR="R5jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"RR&72Qh;R
RRRRRRRRRRMRC8VRH;R
RRRRRRMRC8sRbF#OC#S;
CRM8oCCMsCN0Rcz4;R
RR4Rz6:RRRRHV50MFRM8H_osC2CRoMNCs0RC
RRRRRRRRRHRRMC_so=R<Rj5"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jjR7&RQ;h2
MSC8CRoMNCs0zCR4
6;
RRRRz7ma=R<R0Fk_osC58IH04E-RI8FMR0Fj
2;
RRRR_N8sRCo<q=R7;7)
RRRRR--tCCMsCN0RC0ERv)qRDOCDN#RM#8RCODC0FRDoRHOVRFs)Aqv41n_44_1
RRRRUz4RH:RVOR5EOFHCH_I8R0E=2R4RMoCC0sNCR
SREzO	RR:H5VRR8N8s8IH0>ERRR4c2CRoMNCs0RC
RRRRRzRRO:D	RFbsO#C#Rp5BiS2
RRRRRCRLo
HMSRRRRRRRH5VRB'piCMPC0MRN8pRBiRR='24'RC0EMR
SRRRRRRRRRsN8CNo58I8sHE80-84RF0IMFcR42=R<R_N8s5CoNs88I0H8ER-48MFI04FRc
2;SRSRR8CMR;HV
CSSMb8RsCFO#k#RO;D	
RSRCRM8oCCMsCN0REzO	R;
RRRRRzRR4:gRRsVFRHHRM8R5CEb0_lMk_DOCD-#RRR428MFI0jFRRMoCC0sNCR
RR-R-RRQV58N8s8IH0>ERR24cRCMC8FR0RCOsNR0CI0sHCMRCNCLDR8NMR0FkbRk0CLMND#CRCODC0FRDo
HORRRRRRRRSjz.RH:RVNR58I8sHE80R4>Rco2RCsMCN
0CSR--VRHGVRFsODNDRU4dUR(,#CCDOF0RVsR0HN#00MCRFL0RCoHMRosCHC#0s
C8RRRRRRRRRRRRRRRRF_k0CHM52=R<R''4RCIEMNR58osC58N8s8IH04E-RI8FMR0F4Rc2=2RHR#CDCjR''R;
RRRRRRRRRRRRRIRRsC0_M25HRR<=WI RERCM5_N8s5CoNs88I0H8ER-48MFI04FRc=2RRRH2CCD#R''j;R
RRRRRRCRSMo8RCsMCNR0Cz;.j
RRRRR--Q5VRNs88I0H8E=R<R24.RRMFI0sHCMRCNCLDRRFsFbk0kC0RMDNLCCR#D0CORoDFHMORCCC88R
RRRRRRRRRR.Rz4RR:H5VRNs88I0H8E=R<R24cRMoCC0sNCR
RRRRRRRRRRRRRRkRF0M_C5RH2<'=R4
';RRRRRRRRRRRRRRRRI_s0CHM52=R<R;W 
RRRRRRRRRRRR8CMRMoCC0sNC.Rz4R;
R-RR-CRtMNCs00CRE)CRqOvRC#DDR8NMRH0s-N#00
C#RRRRRRRRS.z.RV:RF[sRRRHM58IH0ME_kOl_C#DDR4-R2FR8IFM0RojRCsMCN
0CSNSS0H0sLCk0R_GObbsF#VRFRqA)vn_4dXUc4RR:DCNLD#RHR)"1e=qp"RR&#NsPD+5[4&2RRR",Wa)Q m_v7" =RI&RsF_l8
C;RRRRRRRRRRRRNs00H0LkC3R\s_NlF#VVCR0\FAVR)_qv4UndcRX4:NRDLRCDH"#RA"1aRH&RMo0CCHs'lCNo58IH0RE2&7R""RR&HCM0o'CsHolNC*5H4Undc&2RR""WRH&RMo0CCHs'lCNo5R[2& R""RR&HCM0o'CsHolNCC5o0M_C8C_8b50E5+HRR*424Undc8,RCEb02&2RR""XRH&RMo0CCHs'lCNo54[+2S;
SCSLo
HMRRRRRRRRRRRRSqA)vn_4dXUc4RR:)Aqv41n_4R
SRRRRRRRRRbRRFRs0lRNb557Qj=2R>MRH_osC5,[2R7q7)>R=RIDF_8N8sd54RI8FMR0FjR2, =hR>hR ,1R1)>R=Ra)1,S
SS SWRR=>I_s0CHM52B,Rp=iR>pRBi7,Rm25jRR=>F_k0L4k#5[H,2
2;RRRRRRRRRRRRRRRRF_k0s5Co[<2R=kRF0k_L#H45,R[2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRMSC8CRoMNCs0zCR.
.;RRRRRRRRCRM8oCCMsCN0Rgz4;R
RRMRC8CRoMNCs0zCR4RU;R
RRRRRRRRR
R-RR-CRtMNCs00CRE)CRqOvRC#DDR8NMRD#CCRO0DHFoOFRVsqR)vnA4_
1.Sdz.RH:RVOR5EOFHCH_I8R0E=2R.RMoCC0sNCS
S-V-RHVGRFOsRNRDD4UdU(#,RCODC0VRFRH0s#00NCFRM0CRLHRMosHCo#s0CCS8
RORzE:	RRRHV58RN8HsI8R0E>dR42CRoMNCs0RC
RRRRRzRRO:D	RFbsO#C#Rp5BiS2
RRRRRCRLo
HMSRRRRRRRH5VRB'piCMPC0MRN8pRBiRR='24'RC0EMR
SRRRRRRRRRsN8CNo58I8sHE80-84RF0IMFdR42=R<R_N8s5CoNs88I0H8ER-48MFI04FRd
2;SRSRR8CMR;HV
CSSMb8RsCFO#k#RO;D	
RSRCRM8oCCMsCN0REzO	R;
RSRRzR.c:FRVsRRHH5MR80CbEk_MlC_ODRD#-2R4RI8FMR0FjCRoMNCs0SC
-Q-RVNR58I8sHE80R4>RdM2RCRC80OFRs0CNCsRIHR0CCLMNDNCRMF8Rkk0b0MRCNCLDRD#CCRO0DHFoOR
RRRRRRzRS.:6RRRHV58N8s8IH0>ERR24dRMoCC0sNC-
S-HRVGFRVsNROD4DRd(UU,CR#D0CORRFV0#sH0CN0R0MFRHLCMsoRC#oH0CCs8R
RRRRRRRRRRRRRRkRF0M_C5RH2<'=R4I'RERCM5sN8CNo58I8sHE80-84RF0IMFdR42RR=HC2RDR#C';j'
RRRRRRRRRRRRRRRR0Is_5CMH<2R= RWRCIEMNR58C_so85N8HsI8-0E4FR8IFM0R24dRH=R2DRC#'CRj
';RRRRRRRRS8CMRMoCC0sNC.Rz6S;
-Q-RVNR58I8sHE80RR<=4Rd2MIFRsCH0RNCMLRDCFFsRkk0b0MRCNCLDRD#CCRO0DHFoOCRMC88C
RRSRSRRzR.n:VRHR85N8HsI8R0E<4=Rdo2RCsMCN
0CSRRRRRRRRRRRR0Fk_5CMH<2R=4R''R;
RRRRRRRRRRRRRIRRsC0_M25HRR<=W
 ;RRRRRRRRS8CMRMoCC0sNC.RznS;
-t-RCsMCNR0C0REC)RqvODCD#MRN8sR0H0-#N#0C
RRRRRRRR.Sz(RR:VRFs[MRHRH5I8_0EM_klODCD#RR-482RF0IMFRRjoCCMsCN0
SSSNs00H0LkCORG_FbsbF#RV)RAqUv_4Xg..RR:DCNLD#RHR)"1e=qp"RR&#NsPD*5.[R+.8MFI0.FR*4[+2RR&"W,R) Qa_7vm R="&sRI_8lFCR;
RRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)RAqUv_4Xg..RR:DCNLD#RHR1"Aa&"RR0HMCsoC'NHloIC5HE802RR&"R7"&MRH0CCosl'HN5oCH4*UgR.2&WR""RR&HCM0o'CsHolNC*5[.&2RR"" RH&RMo0CCHs'lCNo50oC_8CM_b8C05E5HRR+4U2*4,g.Rb8C02E2R"&RX&"RR0HMCsoC'NHlo5C5[2+4*;.2
SSSLHCoMR
RRRRRRRRRRARS)_qvU.4gX:.RRv)qA_4n1R.
RRRRRRRRRRRRRRRRRsbF0NRlb7R5Q>R=R_HMs5Co.+*[4FR8IFM0R[.*2q,R7R7)=D>RFNI_858s48.RF0IMF2Rj,hR RR=> Rh,1R1)=)>R1
a,RRRRRRRRRRRRRRRRRRRRRRRRRRRRW= R>sRI0M_C5,H2RiBpRR=>B,piR57m4=2R>kRF0k_L#H.5,[.*+,42R57mj=2R>kRF0k_L#H.5,*R.[;22
RRRRRRRRRRRRRRRR0Fk_osC5[.*2=R<R0Fk_#Lk.,5H.2*[RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_so*5.[2+4RR<=F_k0L.k#5.H,*4[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRSRRCRM8oCCMsCN0R(z.;R
RRSRRCRM8oCCMsCN0Rcz.;R
RRMRC8CRoMNCs0zCR.Rd;RS

RRRR-t-RCsMCNR0C0REC)RqvODCD#MRN8CR#D0CORoDFHVORF)sRq4vAnc_1
.SzURR:H5VROHEFOIC_HE80Rc=R2CRoMNCs0SC
SR--VRHGVRFsODNDRU4dUR(,#CCDOF0RVsR0HN#00MCRFL0RCoHMRosCHC#0s
C8SzRRORE	:VRHR85N8HsI8R0E>.R42CRoMNCs0RC
RRRRRzRRO:D	RFbsO#C#Rp5BiS2
RRRRRCRLo
HMSRRRRRRRH5VRB'piCMPC0MRN8pRBiRR='24'RC0EMR
SRRRRRRRRRsN8CNo58I8sHE80-84RF0IMF.R42=R<R_N8s5CoNs88I0H8ER-48MFI04FR.
2;SRSRR8CMR;HV
CSSMb8RsCFO#k#RO;D	
RSRCRM8oCCMsCN0REzO	R;
RSRRzR.g:FRVsRRHH5MR80CbEk_MlC_ODRD#-2R4RI8FMR0FjCRoMNCs0SC
-Q-RVNR58I8sHE80R4>R.M2RCRC80OFRs0CNCsRIHR0CCLMNDNCRMF8Rkk0b0MRCNCLDRD#CCRO0DHFoOR
RRRRRRzRSd:jRRRHV58N8s8IH0>ERR24.RMoCC0sNC-
S-HRVGFRVsNROD4DRd(UU,CR#D0CORRFV0#sH0CN0R0MFRHLCMsoRC#oH0CCs8R
RRRRRRRRRRRRRRkRF0M_C5RH2<'=R4I'RERCM5sN8CNo58I8sHE80-84RF0IMF.R42RR=HC2RDR#C';j'
RRRRRRRRRRRRRRRR0Is_5CMH<2R= RWRCIEMNR58C_so85N8HsI8-0E4FR8IFM0R24.RH=R2DRC#'CRj
';RRRRRRRRS8CMRMoCC0sNCdRzjS;
-Q-RVNR58I8sHE80RR<=4R.2MIFRsCH0RNCMLRDCFFsRkk0b0MRCNCLDRD#CCRO0DHFoOCRMC88C
RRSRSRRzRd4:VRHR85N8HsI8R0E<4=R.o2RCsMCN
0CSRRRRRRRRRRRR0Fk_5CMH<2R=4R''R;
RRRRRRRRRRRRRIRRsC0_M25HRR<=W
 ;RRRRRRRRS8CMRMoCC0sNCdRz4S;
-t-RCsMCNR0C0REC)RqvODCD#MRN8sR0H0-#N#0C
RRRRRRRRdSz.RR:VRFs[MRHRH5I8_0EM_klODCD#RR-482RF0IMFRRjoCCMsCN0
SSSNs00H0LkCORG_FbsbF#RV)RAqcv_jXgncRR:DCNLD#RHR)"1e=qp"RR&#NsPD*5c[R+c8MFI0cFR*4[+2RR&"W,R) Qa_7vm R="&sRI_8lFCR;
RRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)RAqcv_jXgncRR:DCNLD#RHR1"Aa&"RR0HMCsoC'NHloIC5HE802RR&"R7"&MRH0CCosl'HN5oCHj*cgRn2&WR""RR&HCM0o'CsHolNC*5[c&2RR"" RH&RMo0CCHs'lCNo50oC_8CM_b8C05E5HRR+4c2*j,gnRb8C02E2R"&RX&"RR0HMCsoC'NHlo5C5[2+4*;c2
SSSLHCoMR
RRRRRRRRRRARS)_qvcnjgX:cRRv)qA_4n1Sc
RRRRRRRRRRRRb0FsRblNRQ57RR=>HsM_Cco5*d[+RI8FMR0Fc2*[,7Rq7=)R>FRDI8_N84s54FR8IFM0R,j2RR h= >Rh1,R1=)R>1R)a
,RSSSSW= R>sRI0M_C5,H2RiBpRR=>B,piR57md=2R>kRF0k_L#Hc5,*Rc[2+d,mR75R.2=F>RkL0_k5#cH*,c[2+.,SR
S7SSm254RR=>F_k0Lck#5cH,*4[+27,Rm25jRR=>F_k0Lck#5RH,c2*[2R;
RRRRRRRRRRRRRFRRks0_Cco5*R[2<F=RkL0_k5#cH*,c[I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Coc+*[4<2R=kRF0k_L#Hc5,[c*+R42IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5[c*+R.2<F=RkL0_k5#cH*,c[2+.RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_so*5c[2+dRR<=F_k0Lck#5cH,*d[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRSRRCRM8oCCMsCN0R.zd;R
RRSRRCRM8oCCMsCN0Rgz.;R
RRMRC8CRoMNCs0zCR.
U;
RSRR-R-RMtCC0sNCER0CqR)vCRODRD#NRM8#CCDOD0RFOoHRsVFRv)qA_4n1Sg
zRdd:VRHRE5OFCHO_8IH0=ERRRg2oCCMsCN0
-SS-HRVGFRVsNROD4DRd(UU,CR#D0CORRFV0#sH0CN0R0MFRHLCMsoRC#oH0CCs8R
SREzO	RR:H5VRR8N8s8IH0>ERR244RMoCC0sNCR
RRRRRRORzDR	:bOsFCR##5iBp2R
SRRRRRoLCHSM
RRRRRHRRVBR5pCi'P0CMR8NMRiBpR'=R4R'20MEC
RSRRRRRRRRRNC8so85N8HsI8-0E4FR8IFM0R244RR<=Ns8_CNo58I8sHE80-84RF0IMF4R42S;
SRRRCRM8H
V;SMSC8sRbF#OC#ORkD
	;SCRRMo8RCsMCNR0Cz	OE;R
RRzRSd:cRRsVFRHHRM8R5CEb0_lMk_DOCD-#RRR428MFI0jFRRMoCC0sNC-
S-VRQR85N8HsI8R0E>4R42CRMC08RFsROCCN0RHIs0CCRMDNLCMRN8kRF00bkRNCMLRDC#CCDOD0RFOoH
RRRRRRRRdSz6RR:H5VRNs88I0H8ERR>4R42oCCMsCN0
-S-RGVHRsVFRDONDdR4U,U(RD#CCRO0F0VRs0H#NR0CMRF0LMCHoCRso0H#C8sC
RRRRRRRRRRRRRRRR0Fk_5CMH<2R=4R''ERIC5MRNC8so85N8HsI8-0E4FR8IFM0R244RH=R2DRC#'CRj
';RRRRRRRRRRRRRRRRI_s0CHM52=R<RRW IMECR85N_osC58N8s8IH04E-RI8FMR0F4R42=2RHR#CDCjR''R;
RRRRRSRRCRM8oCCMsCN0R6zd;-
S-VRQR85N8HsI8R0E<4=R4M2RFsRIHR0CCLMNDFCRskRF00bkRNCMLRDC#CCDOD0RFOoHRCMC8
C8RRSRRzRSd:nRRRHV58N8s8IH0<ER=4R42CRoMNCs0SC
RRRRRRRRRRRRF_k0CHM52=R<R''4;R
RRRRRRRRRRRRRRsRI0M_C5RH2<W=R R;
RRRRRSRRCRM8oCCMsCN0Rnzd;-
S-CRtMNCs00CRE)CRqOvRC#DDR8NMRH0s-N#00
C#RRRRRRRRS(zdRV:RF[sRRRHM58IH0ME_kOl_C#DDR4-R2FR8IFM0RojRCsMCN
0CSNSS0H0sLCk0R_GObbsF#VRFRqA)vj_.cUUXRD:RNDLCRRH#"e1)q"p=R#&RsDPN5[g*+8gRF0IMF*Rg[2+4R"&R,)RWQ_a v m7=&"RR_IslCF8;R
RRRRRRRRRR0RN0LsHkR0C\N3slV_FV0#C\VRFRqA)vj_.cUUXRD:RNDLCRRH#"aA1"RR&HCM0o'CsHolNCH5I820ER"&R7&"RR0HMCsoC'NHloHC5*c.jU&2RR""WRH&RMo0CCHs'lCNo5g[*2RR&"R "&MRH0CCosl'HN5oCo_C0C_M880CbEH55R4+R2j*.cRU,80CbER22&XR""RR&HCM0o'CsHolNC[55+*42g
2;SLSSCMoH
RRRRRRRRRRRR)SAq.v_jXcUURR:)Aqv41n_gR
SRRRRRRRRRbRRFRs0lRNb5R7Q=H>RMC_so*5g[R+(8MFI0gFR*,[2R7q7)>R=RIDF_8N8sj54RI8FMR0FjR2, =hR>hR ,1R1)>R=Ra)1,RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRW =I>RsC0_M25H,pRBi>R=RiBp,mR75R(2=F>RkL0_k5#UH*,U[2+(,mR75Rn2=F>RkL0_k5#UH*,U[2+n,RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRR57m6=2R>kRF0k_L#HU5,[U*+,62R57mc=2R>kRF0k_L#HU5,[U*+,c2R57md=2R>kRF0k_L#HU5,[U*+,d2RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRR7.m52>R=R0Fk_#LkU,5HU+*[.R2,74m52>R=R0Fk_#LkU,5HU+*[4R2,7jm52>R=R0Fk_#LkU,5HU2*[,RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRu7Q5Rj2=H>RMC_so*5g[2+U,mR7u25jRR=>bHNs0L$_k5#UH2,[2R;
RRRRRRRRRRRRRFRRks0_Cgo5*R[2<F=RkL0_k5#UH*,U[I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cog+*[4<2R=kRF0k_L#HU5,[U*+R42IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5[g*+R.2<F=RkL0_k5#UH*,U[2+.RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_so*5g[2+dRR<=F_k0LUk#5UH,*d[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cgo5*c[+2=R<R0Fk_#LkU,5HU+*[cI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cog+*[6<2R=kRF0k_L#HU5,[U*+R62IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5[g*+Rn2<F=RkL0_k5#UH*,U[2+nRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_so*5g[2+(RR<=F_k0LUk#5UH,*([+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cgo5*U[+2=R<RsbNH_0$LUk#5[H,2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRSRRCRM8oCCMsCN0R(zd;R
RRSRRCRM8oCCMsCN0Rczd;R
RRMRC8CRoMNCs0zCRd
d;
RSRR-R-RMtCC0sNCER0CqR)vCRODRD#NRM8#CCDOD0RFOoHRsVFRv)qA_4n1
4USUzdRH:RVOR5EOFHCH_I8R0E=UR42CRoMNCs0SC
SR--VRHGVRFsODNDRU4dUR(,#CCDOF0RVsR0HN#00MCRFL0RCoHMRosCHC#0s
C8SzRRORE	:VRHRN5R8I8sHE80R4>RjRR2oCCMsCN0
RRRRRRRRDzO	b:RsCFO#5#RB2pi
RSRRRRRLHCoMR
SRRRRRVRHRp5BiP'CCRM0NRM8BRpi=4R''02RE
CMSRRRRRRRRNRR8osC58N8s8IH04E-RI8FMR0F4Rj2<N=R8C_so85N8HsI8-0E4FR8IFM0R24j;S
SRCRRMH8RVS;
S8CMRFbsO#C#RDkO	S;
RMRC8CRoMNCs0zCRO;E	
RRRRdSzgRR:VRFsHMRHRC58b_0EM_klODCD#RR-482RF0IMFRRjoCCMsCN0
-S-RRQV58N8s8IH0>ERR24jRCMC8FR0RCOsNR0CI0sHCMRCNCLDR8NMR0FkbRk0CLMND#CRCODC0FRDo
HORRRRRRRRSjzcRH:RVNR58I8sHE80R4>Rjo2RCsMCN
0CSR--VRHGVRFsODNDRU4dUR(,#CCDOF0RVsR0HN#00MCRFL0RCoHMRosCHC#0s
C8RRRRRRRRRRRRRRRRF_k0CHM52=R<R''4RCIEMNR58osC58N8s8IH04E-RI8FMR0F4Rj2=2RHR#CDCjR''R;
RRRRRRRRRRRRRIRRsC0_M25HRR<=WI RERCM5_N8s5CoNs88I0H8ER-48MFI04FRj=2RRRH2CCD#R''j;R
RRRRRRCRSMo8RCsMCNR0Cz;cj
-S-RRQV58N8s8IH0<ER=jR42FRMRHIs0CCRMDNLCsRFR0FkbRk0CLMND#CRCODC0FRDoRHOM8CCCR8
SRRRRcSz4RR:H5VRNs88I0H8E=R<R24jRMoCC0sNCR
SRRRRRRRRRFRRkC0_M25HRR<=';4'
RRRRRRRRRRRRRRRR0Is_5CMH<2R= RW;R
RRRRRRCRSMo8RCsMCNR0Cz;c4
-S-RMtCC0sNCER0CqR)vCRODRD#NRM80-sH#00NCR#
RRRRRSRRzRc.:FRVsRR[H5MRI0H8Ek_MlC_ODRD#-2R4RI8FMR0FjCRoMNCs0SC
S0SN0LsHkR0CGbO_s#FbRRFVAv)q_.4jcnX4RD:RNDLCRRH#"e1)q"p=R#&RsDPN5*4U[U+4RI8FMR0F4[U*+R42&,R"RQW)av _m=7 "RR&Ils_F;8C
RRRRRRRRRRRR0N0skHL0\CR3lsN_VFV#\C0RRFVAv)q_.4jcnX4RD:RNDLCRRH#"aA1"RR&HCM0o'CsHolNCH5I820ER"&R7&"RR0HMCsoC'NHloHC5*.4jc&2RR""WRH&RMo0CCHs'lCNo54[*U&2RR"" RH&RMo0CCHs'lCNo50oC_8CM_b8C05E5HRR+442*j,.cRb8C02E2R"&RX&"RR0HMCsoC'NHlo5C5[2+4*24U;S
SSoLCHRM
RRRRRRRRRSRRAv)q_.4jcnX4R):Rq4vAn4_1UR
RRRRRRRRRRRRRRRRRb0FsRblNRQ57RR=>HsM_C4o5U+*[486RF0IMFUR4*,[2R7q7)>R=RIDF_8N8sR5g8MFI0jFR2 ,Rh>R=R, hR)11RR=>),1aRR
RRRRRRRRRRRRRRRRRRRRRRRRRR RWRR=>I_s0CHM52B,Rp=iR>pRBi7,Rm6542>R=R0Fk_#Lk4Hn5,*4n[6+427,Rmc542>R=R0Fk_#Lk4Hn5,*4n[c+42
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRR74m5d=2R>kRF0k_L#54nHn,4*4[+dR2,74m5.=2R>kRF0k_L#54nHn,4*4[+.R2,74m54=2R>kRF0k_L#54nHn,4*4[+4R2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRR57m4Rj2=F>RkL0_kn#454H,n+*[4,j2R57mg=2R>kRF0k_L#54nHn,4*g[+27,Rm25URR=>F_k0L4k#n,5H4[n*+,U2
RRRRRRRRRRRRRRRRRRRRRRRRRRRR57m(=2R>kRF0k_L#54nHn,4*([+27,Rm25nRR=>F_k0L4k#n,5H4[n*+,n2R57m6=2R>kRF0k_L#54nHn,4*6[+2S,
SRSRRmR75Rc2=F>RkL0_kn#454H,n+*[cR2,7dm52>R=R0Fk_#Lk4Hn5,*4n[2+d,mR75R.2=F>RkL0_kn#454H,n+*[.
2,RRRRRRRRRRRRRRRRRRRRRRRRRRRR74m52>R=R0Fk_#Lk4Hn5,*4n[2+4,mR75Rj2=F>RkL0_kn#454H,n2*[,RR
RRRRRRRRRRRRRRRRRRRRRRRRR7RRQ=uR>MRH_osC5*4U[(+4RI8FMR0F4[U*+24n,R
RRRRRRRRRRRRRRRRRRRRRRRRRRmR7u254RR=>bHNs0L$_kn#45.H,*4[+27,Rmju52>R=RsbNH_0$L4k#n,5H.2*[2R;
RRRRRRRRRRRRRFRRks0_C4o5U2*[RR<=F_k0L4k#n,5H4[n*2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_C4o5U+*[4<2R=kRF0k_L#54nHn,4*4[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_C4o5U+*[.<2R=kRF0k_L#54nHn,4*.[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_C4o5U+*[d<2R=kRF0k_L#54nHn,4*d[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_C4o5U+*[c<2R=kRF0k_L#54nHn,4*c[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_C4o5U+*[6<2R=kRF0k_L#54nHn,4*6[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_C4o5U+*[n<2R=kRF0k_L#54nHn,4*n[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_C4o5U+*[(<2R=kRF0k_L#54nHn,4*([+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_C4o5U+*[U<2R=kRF0k_L#54nHn,4*U[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_C4o5U+*[g<2R=kRF0k_L#54nHn,4*g[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_C4o5U+*[4Rj2<F=RkL0_kn#454H,n+*[4Rj2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*4U[4+42=R<R0Fk_#Lk4Hn5,*4n[4+42ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_C4o5U+*[4R.2<F=RkL0_kn#454H,n+*[4R.2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*4U[d+42=R<R0Fk_#Lk4Hn5,*4n[d+42ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_C4o5U+*[4Rc2<F=RkL0_kn#454H,n+*[4Rc2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*4U[6+42=R<R0Fk_#Lk4Hn5,*4n[6+42ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_C4o5U+*[4Rn2<b=RN0sH$k_L#54nH*,.[I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co4[U*+24(RR<=bHNs0L$_kn#45.H,*4[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRSRRCRM8oCCMsCN0R.zc;R
RRSRRCRM8oCCMsCN0Rgzd;R
RRMRC8CRoMNCs0zCRd
U;
RSRR-R-RMtCC0sNCER0CqR)vCRODRD#NRM8#CCDOD0RFOoHRsVFRv)qA_4n1
dnSdzcRH:RVOR5EOFHCH_I8R0E=nRd2CRoMNCs0SC
SR--VRHGVRFsODNDRU4dUR(,#CCDOF0RVsR0HN#00MCRFL0RCoHMRosCHC#0s
C8SzRRORE	:VRHRN5R8I8sHE80Rg>RRo2RCsMCN
0CSRRRRDzO	b:RsCFO#5#RB2pi
RSSRoLCHSM
SRRRH5VRB'piCMPC0MRN8pRBiRR='24'RC0EMS
SRRRRR8RNs5CoNs88I0H8ER-48MFI0gFR2=R<R_N8s5CoNs88I0H8ER-48MFI0gFR2S;
SRRRCRM8H
V;SMSC8sRbF#OC#ORkD
	;SCRRMo8RCsMCNR0Cz	OE;R
SRzRRc:cRRsVFRHHRM8R5CEb0_lMk_DOCD-#RRR428MFI0jFRRMoCC0sNC-
S-VRQR85N8HsI8R0E>2RgRCMC8FR0RCOsNR0CI0sHCMRCNCLDR8NMR0FkbRk0CLMND#CRCODC0FRDo
HOSzSSc:6RRRHV58N8s8IH0>ERRRg2oCCMsCN0
-S-RGVHRsVFRDONDdR4U,U(RD#CCRO0F0VRs0H#NR0CMRF0LMCHoCRso0H#C8sC
SSSS0Fk_5CMH<2R=4R''ERIC5MRNC8so85N8HsI8-0E4FR8IFM0RRg2=2RHR#CDCjR''S;
SISSsC0_M25HRR<=WI RERCM5_N8s5CoNs88I0H8ER-48MFI0gFR2RR=HC2RDR#C';j'
SSSCRM8oCCMsCN0R6zc;-
S-VRQR85N8HsI8R0E<g=R2FRMRHIs0CCRMDNLCsRFR0FkbRk0CLMND#CRCODC0FRDoRHOM8CCCS8
ScSznRR:H5VRNs88I0H8E=R<RRg2oCCMsCN0
SSSS0Fk_5CMH<2R=4R''S;
SISSsC0_M25HRR<=W
 ;SCSSMo8RCsMCNR0Cz;cn
-S-RMtCC0sNCER0CqR)vCRODRD#NRM80-sH#00NCS#
ScSz(RR:VRFs[MRHRH5I8_0EM_klODCD#RR-482RF0IMFRRjoCCMsCN0
SSSNs00H0LkCORG_FbsbF#RV)RAq6v_4d.X.RR:DCNLD#RHR)"1e=qp"RR&#NsPDn5d*d[+nFR8IFM0R*dn[2+4R"&R,)RWQ_a v m7=&"RR_IslCF8;R
RRRRRRRRRR0RN0LsHkR0C\N3slV_FV0#C\VRFRqA)v4_6..XdRD:RNDLCRRH#"aA1"RR&HCM0o'CsHolNCH5I820ER"&R7&"RR0HMCsoC'NHloHC5*.642RR&"RW"&MRH0CCosl'HN5oC[n*d2RR&"R "&MRH0CCosl'HN5oCo_C0C_M880CbEH55R4+R24*6.8,RCEb02&2RR""XRH&RMo0CCHs'lCNo5+5[4d2*n
2;SLSSCMoH
RRRRRRRRRRRRRRRRRRRRRRRRARR)_qv6X4.d:.RRv)qA_4n1
dnRRRRRRRRRRRRRRRRRRRRRRRRRRRRb0FsRblNRQ57RR=>HsM_Cdo5n+*[d84RF0IMFnRd*,[2R7q7)>R=D_FINs8858URF0IMF2Rj,hR RR=> Rh,1R1)=)>R1
a,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR RWRR=>I_s0CHM52B,Rp=iR>pRBi7,Rm45d2>R=R0Fk_#LkdH.5,*d.[4+d27,Rmj5d2>R=R0Fk_#LkdH.5,*d.[j+d2R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR57m.Rg2=F>RkL0_k.#d5dH,.+*[.,g2R57m.RU2=F>RkL0_k.#d5dH,.+*[.,U2R57m.R(2=F>RkL0_k.#d5dH,.+*[.,(2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR7RRmn5.2>R=R0Fk_#LkdH.5,*d.[n+.27,Rm65.2>R=R0Fk_#LkdH.5,*d.[6+.27,Rmc5.2>R=R0Fk_#LkdH.5,*d.[c+.2R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR57m.Rd2=F>RkL0_k.#d5dH,.+*[.,d2R57m.R.2=F>RkL0_k.#d5dH,.+*[.,.2R57m.R42=F>RkL0_k.#d5dH,.+*[.,42
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR7RRmj5.2>R=R0Fk_#LkdH.5,*d.[j+.27,Rmg542>R=R0Fk_#LkdH.5,*d.[g+427,RmU542>R=R0Fk_#LkdH.5,*d.[U+42R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR57m4R(2=F>RkL0_k.#d5dH,.+*[4,(2R57m4Rn2=F>RkL0_k.#d5dH,.+*[4,n2R57m4R62=F>RkL0_k.#d5dH,.+*[4,62
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR7RRmc542>R=R0Fk_#LkdH.5,*d.[c+427,Rmd542>R=R0Fk_#LkdH.5,*d.[d+427,Rm.542>R=R0Fk_#LkdH.5,*d.[.+42
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRmR75244RR=>F_k0Ldk#.,5Hd[.*+244,mR7524jRR=>F_k0Ldk#.,5Hd[.*+24j,mR75Rg2=F>RkL0_k.#d5dH,.+*[gR2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR7RRm25URR=>F_k0Ldk#.,5Hd[.*+,U2R57m(=2R>kRF0k_L#5d.H.,d*([+27,Rm25nRR=>F_k0Ldk#.,5Hd[.*+,n2RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR76m52>R=R0Fk_#LkdH.5,*d.[2+6,mR75Rc2=F>RkL0_k.#d5dH,.+*[cR2,7dm52>R=R0Fk_#LkdH.5,*d.[2+d,RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR57m.=2R>kRF0k_L#5d.H.,d*.[+27,Rm254RR=>F_k0Ldk#.,5Hd[.*+,42R57mj=2R>kRF0k_L#5d.H.,d*,[2RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR7RQu=H>RMC_son5d*d[+6FR8IFM0R*dn[.+d2R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRu7m5Rd2=b>RN0sH$k_L#5d.H*,c[2+d,mR7u25.RR=>bHNs0L$_k.#d5cH,*.[+2R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRu7m5R42=b>RN0sH$k_L#5d.H*,c[2+4,mR7u25jRR=>bHNs0L$_k.#d5cH,*2[2;R
RRRRRRRRRRRRRRRRRRRRRRRRRF_k0s5Cod[n*2=R<R0Fk_#LkdH.5,*d.[I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRRRRRRRRRkRF0C_son5d*4[+2=R<R0Fk_#LkdH.5,*d.[2+4RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRRRRRRRRRF_k0s5Cod[n*+R.2<F=RkL0_k.#d5dH,.+*[.I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRRRRRRRRRkRF0C_son5d*d[+2=R<R0Fk_#LkdH.5,*d.[2+dRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRRRRRRRRRF_k0s5Cod[n*+Rc2<F=RkL0_k.#d5dH,.+*[cI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRRRRRRRRRkRF0C_son5d*6[+2=R<R0Fk_#LkdH.5,*d.[2+6RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRRRRRRRRRF_k0s5Cod[n*+Rn2<F=RkL0_k.#d5dH,.+*[nI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRRRRRRRRRkRF0C_son5d*([+2=R<R0Fk_#LkdH.5,*d.[2+(RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRRRRRRRRRF_k0s5Cod[n*+RU2<F=RkL0_k.#d5dH,.+*[UI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRRRRRRRRRkRF0C_son5d*g[+2=R<R0Fk_#LkdH.5,*d.[2+gRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRRRRRRRRRF_k0s5Cod[n*+24jRR<=F_k0Ldk#.,5Hd[.*+24jRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRRRRRRRRRF_k0s5Cod[n*+244RR<=F_k0Ldk#.,5Hd[.*+244RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRRRRRRRRRF_k0s5Cod[n*+24.RR<=F_k0Ldk#.,5Hd[.*+24.RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRRRRRRRRRF_k0s5Cod[n*+24dRR<=F_k0Ldk#.,5Hd[.*+24dRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRRRRRRRRRF_k0s5Cod[n*+24cRR<=F_k0Ldk#.,5Hd[.*+24cRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRRRRRRRRRF_k0s5Cod[n*+246RR<=F_k0Ldk#.,5Hd[.*+246RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRRRRRRRRRF_k0s5Cod[n*+24nRR<=F_k0Ldk#.,5Hd[.*+24nRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRRRRRRRRRF_k0s5Cod[n*+24(RR<=F_k0Ldk#.,5Hd[.*+24(RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRRRRRRRRRF_k0s5Cod[n*+24URR<=F_k0Ldk#.,5Hd[.*+24URCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRRRRRRRRRF_k0s5Cod[n*+24gRR<=F_k0Ldk#.,5Hd[.*+24gRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRRRRRRRRRF_k0s5Cod[n*+2.jRR<=F_k0Ldk#.,5Hd[.*+2.jRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRRRRRRRRRF_k0s5Cod[n*+2.4RR<=F_k0Ldk#.,5Hd[.*+2.4RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRRRRRRRRRF_k0s5Cod[n*+2..RR<=F_k0Ldk#.,5Hd[.*+2..RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRRRRRRRRRF_k0s5Cod[n*+2.dRR<=F_k0Ldk#.,5Hd[.*+2.dRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRRRRRRRRRF_k0s5Cod[n*+2.cRR<=F_k0Ldk#.,5Hd[.*+2.cRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRRRRRRRRRF_k0s5Cod[n*+2.6RR<=F_k0Ldk#.,5Hd[.*+2.6RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRRRRRRRRRF_k0s5Cod[n*+2.nRR<=F_k0Ldk#.,5Hd[.*+2.nRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRRRRRRRRRF_k0s5Cod[n*+2.(RR<=F_k0Ldk#.,5Hd[.*+2.(RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRRRRRRRRRF_k0s5Cod[n*+2.URR<=F_k0Ldk#.,5Hd[.*+2.URCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRRRRRRRRRF_k0s5Cod[n*+2.gRR<=F_k0Ldk#.,5Hd[.*+2.gRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRRRRRRRRRF_k0s5Cod[n*+2djRR<=F_k0Ldk#.,5Hd[.*+2djRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRRRRRRRRRF_k0s5Cod[n*+2d4RR<=F_k0Ldk#.,5Hd[.*+2d4RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRRRRRRRRRF_k0s5Cod[n*+2d.RR<=bHNs0L$_k.#d5cH,*R[2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[dRd2<b=RN0sH$k_L#5d.H*,c[2+4RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRRRRRRRRRF_k0s5Cod[n*+2dcRR<=bHNs0L$_k.#d5cH,*.[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRRRRRRRRR0Fk_osC5*dn[6+d2=R<RsbNH_0$Ldk#.,5Hc+*[dI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';SCSSMo8RCsMCNR0Cz;c(
CSSMo8RCsMCNR0Cz;cc
MSC8CRoMNCs0zCRc
d;
8CMRONsECH0Os0kCDRLF_O	s;Nl
s
NO0EHCkO0sMCRFI_s_COEOF	RVqR)v)h_W#RH
MVkOF0HMkRVMHO_M5H0LRR:LDFFC2NMR0sCkRsM#H0sMHoR#C
Lo
HMRVRHR25LRC0EMR
RRCRs0Mks5F"hRNsC8s/IHR0COVFMD0HORCOEOR	31kHlDHN0FlMRHN#l0ROEb#F#HCLDR"!!2R;
R#CDCR
RRCRs0Mks5M"'FI_s_COEOR	'H0#RE#CRNRlCN'#RLODF	N_slV'RF#sRHDMoCFRbs)0Rq"v#2R;
R8CMR;HV
8CMRMVkOM_HH
0;Ns00H0LkCCRoMNCs0_FssFCbs:0RRs#0H;Mo
N--0H0sLCk0RMoCC0sNFss_CsbF0VRFR_MFsOI_E	CORN:RsHOE00COkRsCHV#Rk_MOH0MH58N8sC_so
2;VOkM0MHFRs#0H.Mo#5DPNRR:#H0sMRo2skC0s#MR0D8_FOoH_OPC0RFsHP#
NNsHLRDC#RDP:0R#8F_Do_HOP0COFNs5'oEHE'-NDRFI8MFI0jFR2P;
NNsHLRDCHRR:HCM0o;Cs
oLCHRM
RsVFRHHRMRRj0#FRDEP'HRoEDbFF
RRRRRHV5NN5'oEHE2-HR'=R4R'20MEC
RSR#5DPH:2R=4R''S;
CCD#
RSR#5DPH:2R=jR''S;
CRM8H
V;RMRC8FRDF
b;RCRs0MksRP#D;M
C80R#soHM.P#D;k
VMHO0F#MRD#P.0MsHoR5N:0R#8F_Do_HOP0COFRs2skC0s#MR0MsHo#RH
sPNHDNLCRR#:0R#soHM5EN'H-oENF'DIR+48MFI04FR2P;
NNsHLRDCHRR:HCM0o;Cs
oLCHRM
RsVFRHHRM'RNDRFI0NFR'oEHEFRDFRb
RHRRVNR55RH2=4R''02RE
CMS#RR5NH-'IDF+R42:'=R4
';S#CDCR
SRH#5-DN'F4I+2=R:R''j;C
SMH8RVR;
R8CMRFDFbR;
R0sCkRsM#C;
M#8RD#P.0MsHoN;
0H0sLCk0R_GObbsF#RR:#H0sM
o;-F-OMN#0M#0RsDPNR#:R0D8_FOoH_OPC05FsI0H8ER-48MFI0jFR2=R:Rs#0H.Mo#5DPs_#08NN02-;
-CRLoRHMLODF	NRsllRHblDCCNM00MHFRo#HM#ND
MVkOF0HMCRo0E_OFCHO_8IH0IE5HE80RH:RMo0CCRs2skC0sHMRMo0CCHsR#N
PsLHNDPCRN:DRR0HMCsoCRR:=jP;
NNsHLRDC8dHP.8,RHnP4,HR8PRU,8cHP,HR8PR.,84HPRH:RMo0CC
s;LHCoMR
R8dHP.=R:RH5I8-0E4d2/nR;
RP8H4:nR=IR5HE80-/424
U;RHR8P:UR=IR5HE80-/42gR;
RP8Hc=R:RH5I8-0E4c2/;R
R8.HPRR:=58IH04E-2;/.
8RRHRP4:5=RI0H8E2-4;R
RH5VR84HPRj>R2ER0CRM
RPRRN:DR=NRPDRR+4R;
R8CMR;HV
HRRV8R5HRP.>2RjRC0EMR
RRNRPD=R:RDPNR4+R;R
RCRM8H
V;RVRHRH58P>cRRRj20MEC
RRRRDPNRR:=PRND+;R4
CRRMH8RVR;
RRHV5P8HURR>j02RE
CMRRRRPRND:P=RN+DRR
4;RMRC8VRH;R
RH5VR84HPnRR>j02RE
CMRRRRPRND:P=RN+DRR
4;RMRC8VRH;-
-RVRHRH58PRd.>2RjRC0EM-
-RRRRPRND:P=RN+DRR
4;-R-RCRM8H
V;RVRHRN5PDRR>.02RERCM
RRRR0sCkRsM5*.R*NRPDRR+.*R*RN5PDRR-d;22
CRRD
#CRRRRskC0s5MR.*R*RDPN2R;
R8CMR;HV
8CMR0oC_FOEH_OCI0H8EV;
k0MOHRFMo_C0OHEFO8C_CEb05b8C0:ERR0HMCsoC2CRs0MksR0HMCsoCR
H#PHNsNCLDRO8_EOFHCC_8bR0E:MRH0CCos=R:R
j;LHCoMR
RH5VR80CbERR>U.4g2ER0CRM
R8RR_FOEH_OC80CbE=R:Rd4nU
c;RDRC#RHV5b8C0<ER=4RUgN.RM88RCEb0Rc>RjRgn2ER0CRM
R8RR_FOEH_OC80CbE=R:RgU4.R;
R#CDH5VR80CbE=R<RgcjnMRN8CR8bR0E>jR.cRU20MEC
RRRRO8_EOFHCC_8bR0E:c=Rj;gn
CRRDV#HRC58bR0E<.=RjRcUNRM880CbERR>4cj.R02RE
CMRRRR8E_OFCHO_b8C0:ER=jR.c
U;RDRC#RHV5b8C0<ER=jR4.NcRM88RCEb0R6>R4R.20MEC
RRRRO8_EOFHCC_8bR0E:4=Rj;.c
CRRDV#HRC58bR0E<6=R4R.20MEC
RRRRO8_EOFHCC_8bR0E:6=R4
.;RMRC8VRH;R
RskC0s8MR_FOEH_OC80CbEC;
Mo8RCO0_EOFHCC_8b;0E
MVkOF0HMCRo0H_I8_0El_F8UE5OFCHO_RI8:MRH0CCoss2RCs0kMMRH0CCos#RH
sPNHDNLCHRI8_0El_F8URR:HCM0o;Cs
oLCHRM
RRHV5FOEH_OCI>8RRRU20MEC
RRRR8IH0lE_FU8_RR:=OHEFOIC_8RR-5FOEH_OCIl8RFU8R2R;
R#CDCR
RRHRI8_0El_F8U=R:RFOEH_OCI
8;RMRC8VRH;R
RskC0sIMRHE80_8lF_
U;CRM8o_C0I0H8EF_l8;_U
F
OMN#0MI0R_FOEH_OCI0H8ERR:HCM0oRCs:o=RCO0_EOFHCH_I850EI0H8E
2;O#FM00NMROI_EOFHCC_8bR0E:MRH0CCos=R:Rd4nUoc/CI0_HE80_8lF_IU5_FOEH_OCI0H8E
2;O#FM00NMRO8_EOFHCC_8bR0E:MRH0CCos=R:R0oC_FOEH_OC80CbEC58b20E;F
OMN#0M80R_FOEH_OCI0H8ERR:HCM0oRCs:5=R4Undc_/8OHEFO8C_CEb02RR+5n54d/Uc8E_OFCHO_b8C0RE2/2RU;V

k0MOHRFMo_C0M_klODCD#85IRH:RMo0CCOs;EOFHC8_IRH:RMo0CCRs2skC0sHMRMo0CCHsR#N
PsLHNDMCRkOl_C#DDRH:RMo0CC
s;LHCoMR
RM_klODCD#=R:R85I-/42OHEFOIC_8RR+4R;
R0sCkRsMM_klODCD#C;
Mo8RCM0_kOl_C#DD;V

k0MOHRFMo_C0#CHx5OIMRH:RMo0CCRs;8RMO:MRH0CCoss2RCs0kMMRH0CCos#RH
oLCHRM
RCRs0MksROIMR8*RM
O;CRM8o_C0#CHx;V

k0MOHRFMo_C0LDFF8_58#CHxRH:RMo0CCRs;IH_#x:CRR0HMCsoC;_R8O:IRR0HMCsoC;_RIO:IRR0HMCsoC2CRs0MksR0HMCsoCR
H#LHCoMV
HR_58#CHxRR<=IH_#xRC20MEC
sRRCs0kM_R8O
I;CCD#
sRRCs0kM_RIO
I;CRM8H
V;CRM8o_C0LDFF8V;
k0MOHRFMo_C0C_M880CbEH5#x:CRR0HMCsoCR8;RCEb0RH:RMo0CCRs2skC0sHMRMo0CCHsR#N
PsLHNDlCRH#M_HRxC:MRH0CCos=R:R
j;LHCoMR
Rl_HM#CHxRR:=80CbER;
RRHV5x#HCRR<80CbE02RE
CMRRRRl_HM#CHxRR:=#CHx;R
RCRM8H
V;RCRs0MksRMlH_x#HCC;
Mo8RCC0_M88_CEb0;O

F0M#NRM0OHEFOIC_HE80RH:RMo0CC:sR=CRo0F_LF5D8o_C0#CHx50oC_lMk_DOCDI#5HE80,_R8OHEFOIC_HE802C,o0k_MlC_OD5D#80CbE8,R_FOEH_OC80CbE,22
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRCRo0H_#xoC5CM0_kOl_C#DD58IH0RE,IE_OFCHO_8IH0,E2o_C0M_klODCD#C58b,0EROI_EOFHCC_8b20E2S,
SSSSSSSSS8SR_FOEH_OCI0H8EI,R_FOEH_OCI0H8E
2;O#FM00NMR8IH0ME_kOl_C#DDRH:RMo0CC:sR=CRo0F_LF5D8o_C0#CHx50oC_lMk_DOCDI#5HE80,_R8OHEFOIC_HE802C,o0k_MlC_OD5D#80CbE8,R_FOEH_OC80CbE,22
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR0oC_x#HCC5o0k_MlC_OD5D#I0H8EI,R_FOEH_OCI0H8Eo2,CM0_kOl_C#DD5b8C0RE,IE_OFCHO_b8C02E2,S
SSSSSSSSSSRRRRH5I8-0E482/_FOEH_OCI0H8E5,RI0H8E2-4/OI_EOFHCH_I820ER4+R;F
OMN#0M80RCEb0_lMk_DOCD:#RR0HMCsoCRR:=o_C0LDFF8C5o0H_#xoC5CM0_kOl_C#DD58IH0RE,8E_OFCHO_8IH0,E2o_C0M_klODCD#C58b,0ERO8_EOFHCC_8b20E2R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRCRo0H_#xoC5CM0_kOl_C#DD58IH0RE,IE_OFCHO_8IH0,E2o_C0M_klODCD#C58b,0EROI_EOFHCC_8b20E2S,
SSSSSSSSSRRR5b8C04E-2_/8OHEFO8C_CEb0,8R5CEb0-/42IE_OFCHO_b8C0RE2+;R4SOR
F0M#NRM0xFCsR#:R0D8_FOoH_OPC05FsOHEFOIC_HE80*8IH0ME_kOl_C#DD-8IH04E-RI8FMR0Fj:2R=FR50sEC#>R=R''j2O;
F0M#NRM0#NsPDD_#PRR:#_08DHFoOC_POs0F5FOEH_OCI0H8EH*I8_0EM_klODCD#R-48MFI0jFR2=R:RsxCFRR&#H0sM#o.DsP5#80_N20N;F
OMN#0M#0RsDPNR#:R0MsHoE5OFCHO_8IH0IE*HE80_lMk_DOCD8#RF0IMF2R4RR:=#.DP#H0sM#o5sDPN_P#D2-;
-o#HM#NDRsVFRMMF-ED#N8bCRFLDOs	RN
l#0C$bR0Fk_#Lk4$_0bHCR#sRNsRN$5b8C0ME_kOl_C#DD-84RF0IMF,RjR8IH0ME_kOl_C#DD-84RF0IMF2RjRRFV#_08DHFoO#;
HNoMDkRF0k_L#:4RR0Fk_#Lk4$_0bRC;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-7R.RsNsNF$RVFR8k50RHkMb0FR0RH0s-N#002C#
b0$CkRF0k_L#0._$RbCHN#Rs$sNRC58b_0EM_klODCD#R-48MFI0jFR,*R.I0H8Ek_MlC_OD+D#4FR8IFM0RRj2F#VR0D8_FOoH;H
#oDMNR0Fk_#Lk.RR:F_k0L.k#_b0$CR;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RR.7NNss$VRFRk8F0HR5M0bkRR0F0-sH#00NC
#20C$bR0Fk_#Lkc$_0bHCR#sRNsRN$5b8C0ME_kOl_C#DD-84RF0IMF,RjRIc*HE80_lMk_DOCDd#+RI8FMR0FjF2RV0R#8F_Do;HO
o#HMRNDF_k0Lck#RF:RkL0_k_#c0C$b;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--.N7Rs$sNRRFV80FkRM5HbRk000FRs#H-0CN0#02
$RbCF_k0LUk#_b0$C#RHRsNsN5$R80CbEk_MlC_OD-D#4FR8IFM0RRj,UH*I8_0EM_klODCD#R+(8MFI0jFR2VRFR8#0_oDFH
O;#MHoNFDRkL0_kR#U:kRF0k_L#0U_$;bCRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-.-R7sRNsRN$F8VRFRk05bHMk00RFsR0H0-#N#0C2$
0bbCRN0sH$k_L#0U_$RbCHN#Rs$sNRC58b_0EM_klODCD#R-48MFI0jFR,HRI8_0EM_klODCD#R-48MFI0jFR2VRFR8#0_oDFH
O;#MHoNbDRN0sH$k_L#:URRsbNH_0$LUk#_b0$CR;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-.-R7sRNsRN$F8VRFRk05bHMk00RFsR0H0-#N#0C2$
0bFCRkL0_kn#4_b0$C#RHRsNsN5$R80CbEk_MlC_OD-D#4FR8IFM0RRj,4In*HE80_lMk_DOCD4#+6FR8IFM0RRj2F#VR0D8_FOoH;H
#oDMNR0Fk_#Lk4:nRR0Fk_#Lk40n_$;bCRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-.-R7sRNsRN$F8VRFRk05bHMk00RFsR0H0-#N#0C2$
0bbCRN0sH$k_L#_4n0C$bRRH#NNss$8R5CEb0_lMk_DOCD4#-RI8FMR0Fj.,R*8IH0ME_kOl_C#DD+84RF0IMF2RjRRFV#_08DHFoO#;
HNoMDNRbs$H0_#Lk4:nRRsbNH_0$L4k#n$_0bRC;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-7R.RsNsNF$RVFR8k50RHkMb0FR0RH0s-N#002C#
b0$CkRF0k_L#_d.0C$bRRH#NNss$8R5CEb0_lMk_DOCD4#-RI8FMR0Fjd,R.H*I8_0EM_klODCD#4+dRI8FMR0FjF2RV0R#8F_Do;HO
o#HMRNDF_k0Ldk#.RR:F_k0Ldk#.$_0bRC;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-7R.RsNsNF$RVFR8k50RHkMb0FR0RH0s-N#002C#
b0$CNRbs$H0_#Lkd0._$RbCHN#Rs$sNRC58b_0EM_klODCD#R-48MFI0jFR,*RcI0H8Ek_MlC_OD+D#dFR8IFM0RRj2F#VR0D8_FOoH;H
#oDMNRsbNH_0$Ldk#.RR:bHNs0L$_k.#d_b0$CR;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RR.7NNss$VRFRk8F0HR5M0bkRR0F0-sH#00NC
#2#MHoNFDRkC0_MRR:#_08DHFoOC_POs0F5b8C0ME_kOl_C#DD-84RF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RNCML#DCRsVFRH0s-N#00
C##MHoNIDRsC0_MRR:#_08DHFoOC_POs0F5b8C0ME_kOl_C#DD-84RF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RHIs0CCRMDNLCV#RFCsRNROEsRFIF)VRqOvRC#DD
o#HMRNDHsM_C:oRR8#0_oDFHPO_CFO0sH5I8+0Ed86RF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-k-R#RC80sFRC#oH0RCs7RQh
o#HMRNDF_k0sRCo:0R#8F_Do_HOP0COFIs5HE80+Rd68MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-k-R#RC80sFRC#oH0RCs7amz
o#HMRNDNs8_C:oRR8#0_oDFHPO_CFO0s85N8HsI8-0E4FR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-#RkC08RFCRso0H#CqsR7
7)#MHoNDDRFNI_8R8s:0R#8F_Do_HOP0COF4s5dFR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-8RN8LsRHR0#HkMb0FR0Rv)qRDOCD5#RcHRL0s#RCHJks2C8
o#HMRNDNC8soRR:#_08DHFoOC_POs0F58N8s8IH04E-RI8FMR0FjR2;-0-RFCRso0H#C0sRE#CRCODC0HR#oDMNRRFV0#sH0CN0
R--CRM8LODF	NRsllRHblDCCNM00MHFRo#HM#ND
0N0skHL0\CR3lsN_VFV#\C0R#:R0MsHo
;
LHCoMR
R
RRRRR--QNVR8I8sHE80RO<REOFHCH_I8R0ENH##o'MRj0'RFMRkk8#CR0LH#R
RRjRzRRR:H5VRNs88I0H8ERR=4o2RCsMCN
0CSRRRRIDF_8N8s=R<Rj"jjjjjjjjjj"jjRN&R8C_so25j;C
SMo8RCsMCNR0Cz
j;RRRRzR4R:VRHR85N8HsI8R0E=2R.RMoCC0sNCR
SRDRRFNI_8R8s<"=Rjjjjjjjjjjjj"RR&Ns8_C4o5RI8FMR0Fj
2;S8CMRMoCC0sNC4Rz;R
RR.RzRRR:H5VRNs88I0H8ERR=do2RCsMCN
0CSRRRRIDF_8N8s=R<Rj"jjjjjjjjjj&"RR_N8s5Co.FR8IFM0R;j2
MSC8CRoMNCs0zCR.R;
RzRRd:RRRRHV58N8s8IH0=ERRRc2oCCMsCN0
RSRRFRDI8_N8<sR=jR"jjjjjjjjj&"RR_N8s5CodFR8IFM0R;j2
MSC8CRoMNCs0zCRdR;
RzRRc:RRRRHV58N8s8IH0=ERRR62oCCMsCN0
RSRRFRDI8_N8<sR=jR"jjjjjjjj"RR&Ns8_Cco5RI8FMR0Fj
2;S8CMRMoCC0sNCcRz;R
RR6RzRRR:H5VRNs88I0H8ERR=no2RCsMCN
0CSRRRRIDF_8N8s=R<Rj"jjjjjjRj"&8RN_osC586RF0IMF2Rj;C
SMo8RCsMCNR0Cz
6;RRRRzRnR:VRHR85N8HsI8R0E=2R(RMoCC0sNCR
SRDRRFNI_8R8s<"=Rjjjjj"jjRN&R8C_soR5n8MFI0jFR2S;
CRM8oCCMsCN0R;zn
RRRRRz(RH:RVNR58I8sHE80RU=R2CRoMNCs0SC
RRRRD_FINs88RR<="jjjj"jjRN&R8C_soR5(8MFI0jFR2S;
CRM8oCCMsCN0R;z(
RRRRRzURH:RVNR58I8sHE80Rg=R2CRoMNCs0SC
RRRRD_FINs88RR<="jjjjRj"&8RN_osC58URF0IMF2Rj;C
SMo8RCsMCNR0Cz
U;RRRRzRgR:VRHR85N8HsI8R0E=jR42CRoMNCs0SC
RRRRD_FINs88RR<="jjjj&"RR_N8s5CogFR8IFM0R;j2
MSC8CRoMNCs0zCRgR;
RzRR4RjR:VRHR85N8HsI8R0E=4R42CRoMNCs0SC
RRRRD_FINs88RR<="jjj"RR&Ns8_C4o5jFR8IFM0R;j2
MSC8CRoMNCs0zCR4
j;RRRRzR44RH:RVNR58I8sHE80R4=R.o2RCsMCN
0CSRRRRIDF_8N8s=R<Rj"j"RR&Ns8_C4o54FR8IFM0R;j2
MSC8CRoMNCs0zCR4
4;RRRRzR4.RH:RVNR58I8sHE80R4=Rdo2RCsMCN
0CSRRRRIDF_8N8s=R<R''jRN&R8C_so.54RI8FMR0Fj
2;S8CMRMoCC0sNC4Rz.R;
RzRR4RdR:VRHR85N8HsI8R0E>dR42CRoMNCs0SC
RRRRD_FINs88RR<=Ns8_C4o5dFR8IFM0R;j2
MSC8CRoMNCs0zCR4
d;
RRRRR--Q5VR8_HMs2CoRosCHC#0sQR7h#RkHRMoB
piRRRRzR4cRH:RV8R5HsM_CRo2oCCMsCN0
RRRRRRRRFbsO#C#Rp5Bi7,RQRh2LHCoMR
RRRRRRRRRRVRHRp5BiRR='R4'NRM8B'piCMPC002RE
CMRRRRRRRRRRRRRRRRHsM_C<oR="R5jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"RR&72Qh;R
RRRRRRRRRRMRC8VRH;R
RRRRRRMRC8sRbF#OC#S;
CRM8oCCMsCN0Rcz4;R
RR4Rz6:RRRRHV50MFRM8H_osC2CRoMNCs0RC
RRRRRRRRRHRRMC_so=R<Rj5"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jjR7&RQ;h2
MSC8CRoMNCs0zCR4
6;
RRRRz7ma=R<R0Fk_osC58IH04E-RI8FMR0Fj
2;
RRRR_N8sRCo<q=R7;7)
RRRRR--tCCMsCN0RC0ERv)qRDOCDN#RM#8RCODC0FRDoRHOVRFs)Aqv41n_44_1
RRRRUz4RH:RVOR5EOFHCH_I8R0E=2R4RMoCC0sNCR
SREzO	RR:H5VRR8N8s8IH0>ERRR4c2CRoMNCs0RC
RRRRRzRRO:D	RFbsO#C#Rp5BiS2
RRRRRCRLo
HMSRRRRRRRH5VRB'piCMPC0MRN8pRBiRR='24'RC0EMR
SRRRRRRRRRsN8CNo58I8sHE80-84RF0IMFcR42=R<R_N8s5CoNs88I0H8ER-48MFI04FRc
2;SRSRR8CMR;HV
CSSMb8RsCFO#k#RO;D	
RSRCRM8oCCMsCN0REzO	R;
RRRRRzRR4:gRRsVFRHHRM8R5CEb0_lMk_DOCD-#RRR428MFI0jFRRMoCC0sNCR
RR-R-RRQV58N8s8IH0>ERR24cRCMC8FR0RCOsNR0CI0sHCMRCNCLDR8NMR0FkbRk0CLMND#CRCODC0FRDo
HORRRRRRRRSjz.RH:RVNR58I8sHE80R4>Rco2RCsMCN
0CSR--VRHGVRFsODNDRU4dUR(,#CCDOF0RVsR0HN#00MCRFL0RCoHMRosCHC#0s
C8RRRRRRRRRRRRRRRRF_k0CHM52=R<R''4RCIEMNR58osC58N8s8IH04E-RI8FMR0F4Rc2=2RHR#CDCjR''R;
RRRRRRRRRRRRRIRRsC0_M25HRR<=WI RERCM5_N8s5CoNs88I0H8ER-48MFI04FRc=2RRRH2CCD#R''j;R
RRRRRRCRSMo8RCsMCNR0Cz;.j
RRRRR--Q5VRNs88I0H8E=R<R24.RRMFI0sHCMRCNCLDRRFsFbk0kC0RMDNLCCR#D0CORoDFHMORCCC88R
RRRRRRRRRR.Rz4RR:H5VRNs88I0H8E=R<R24cRMoCC0sNCR
RRRRRRRRRRRRRRkRF0M_C5RH2<'=R4
';RRRRRRRRRRRRRRRRI_s0CHM52=R<R;W 
RRRRRRRRRRRR8CMRMoCC0sNC.Rz4R;
R-RR-CRtMNCs00CRE)CRqOvRC#DDR8NMRH0s-N#00
C#RRRRRRRRS.z.RV:RF[sRRRHM58IH0ME_kOl_C#DDR4-R2FR8IFM0RojRCsMCN
0CSNSS0H0sLCk0R_GObbsF#VRFRqA)vn_4dXUc4RR:DCNLD#RHR)"1e=qp"RR&#NsPD+5[4&2RRR",Wa)Q m_v7" =RI&RsF_l8
C;RRRRRRRRRRRRNs00H0LkC3R\s_NlF#VVCR0\FAVR)_qv4UndcRX4:NRDLRCDH"#RA"1aRH&RMo0CCHs'lCNo58IH0RE2&7R""RR&HCM0o'CsHolNC*5H4Undc&2RR""WRH&RMo0CCHs'lCNo5R[2& R""RR&HCM0o'CsHolNCC5o0M_C8C_8b50E5+HRR*424Undc8,RCEb02&2RR""XRH&RMo0CCHs'lCNo54[+2S;
SCSLo
HMRRRRRRRRRRRRSqA)vn_4dXUc4RR:)Aqv41n_4R
SRRRRRRRRRbRRFRs0lRNb557Qj=2R>MRH_osC5,[2R7q7)>R=RIDF_8N8sd54RI8FMR0FjR2, =hR>hR ,1R1)>R=Ra)1,S
SS SWRR=>I_s0CHM52B,Rp=iR>pRBi7,Rm25jRR=>F_k0L4k#5[H,2
2;RRRRRRRRRRRRRRRRF_k0s5Co[<2R=kRF0k_L#H45,R[2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRMSC8CRoMNCs0zCR.
.;RRRRRRRRCRM8oCCMsCN0Rgz4;R
RRMRC8CRoMNCs0zCR4RU;R
RRRRRRRRR
R-RR-CRtMNCs00CRE)CRqOvRC#DDR8NMRD#CCRO0DHFoOFRVsqR)vnA4_
1.Sdz.RH:RVOR5EOFHCH_I8R0E=2R.RMoCC0sNCS
S-V-RHVGRFOsRNRDD4UdU(#,RCODC0VRFRH0s#00NCFRM0CRLHRMosHCo#s0CCS8
RORzE:	RRRHV58RN8HsI8R0E>dR42CRoMNCs0RC
RRRRRzRRO:D	RFbsO#C#Rp5BiS2
RRRRRCRLo
HMSRRRRRRRH5VRB'piCMPC0MRN8pRBiRR='24'RC0EMR
SRRRRRRRRRsN8CNo58I8sHE80-84RF0IMFdR42=R<R_N8s5CoNs88I0H8ER-48MFI04FRd
2;SRSRR8CMR;HV
CSSMb8RsCFO#k#RO;D	
RSRCRM8oCCMsCN0REzO	R;
RSRRzR.c:FRVsRRHH5MR80CbEk_MlC_ODRD#-2R4RI8FMR0FjCRoMNCs0SC
-Q-RVNR58I8sHE80R4>RdM2RCRC80OFRs0CNCsRIHR0CCLMNDNCRMF8Rkk0b0MRCNCLDRD#CCRO0DHFoOR
RRRRRRzRS.:6RRRHV58N8s8IH0>ERR24dRMoCC0sNC-
S-HRVGFRVsNROD4DRd(UU,CR#D0CORRFV0#sH0CN0R0MFRHLCMsoRC#oH0CCs8R
RRRRRRRRRRRRRRkRF0M_C5RH2<'=R4I'RERCM5sN8CNo58I8sHE80-84RF0IMFdR42RR=HC2RDR#C';j'
RRRRRRRRRRRRRRRR0Is_5CMH<2R= RWRCIEMNR58C_so85N8HsI8-0E4FR8IFM0R24dRH=R2DRC#'CRj
';RRRRRRRRS8CMRMoCC0sNC.Rz6S;
-Q-RVNR58I8sHE80RR<=4Rd2MIFRsCH0RNCMLRDCFFsRkk0b0MRCNCLDRD#CCRO0DHFoOCRMC88C
RRSRSRRzR.n:VRHR85N8HsI8R0E<4=Rdo2RCsMCN
0CSRRRRRRRRRRRR0Fk_5CMH<2R=4R''R;
RRRRRRRRRRRRRIRRsC0_M25HRR<=W
 ;RRRRRRRRS8CMRMoCC0sNC.RznS;
-t-RCsMCNR0C0REC)RqvODCD#MRN8sR0H0-#N#0C
RRRRRRRR.Sz(RR:VRFs[MRHRH5I8_0EM_klODCD#RR-482RF0IMFRRjoCCMsCN0
SSSNs00H0LkCORG_FbsbF#RV)RAqUv_4Xg..RR:DCNLD#RHR)"1e=qp"RR&#NsPD*5.[R+.8MFI0.FR*4[+2RR&"W,R) Qa_7vm R="&sRI_8lFCR;
RRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)RAqUv_4Xg..RR:DCNLD#RHR1"Aa&"RR0HMCsoC'NHloIC5HE802RR&"R7"&MRH0CCosl'HN5oCH4*UgR.2&WR""RR&HCM0o'CsHolNC*5[.&2RR"" RH&RMo0CCHs'lCNo50oC_8CM_b8C05E5HRR+4U2*4,g.Rb8C02E2R"&RX&"RR0HMCsoC'NHlo5C5[2+4*;.2
SSSLHCoMR
RRRRRRRRRRARS)_qvU.4gX:.RRv)qA_4n1S.
RRRRRRRRRRRRb0FsRblNRQ57RR=>HsM_C.o5*4[+RI8FMR0F.2*[,7Rq7=)R>FRDI8_N84s5.FR8IFM0R,j2RR h= >Rh1,R1=)R>1R)aS,
SWSS >R=R0Is_5CMHR2,BRpi=B>RpRi,74m52>R=R0Fk_#Lk.,5H.+*[4R2,7jm52>R=R0Fk_#Lk.,5HR[.*2
2;RRRRRRRRRRRRRRRRF_k0s5Co.2*[RR<=F_k0L.k#5.H,*R[2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5[.*+R42<F=RkL0_k5#.H*,.[2+4RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRCRSMo8RCsMCNR0Cz;.(
RRRRCRSMo8RCsMCNR0Cz;.c
RRRR8CMRMoCC0sNC.RzdR;R
R
SR-RR-CRtMNCs00CRE)CRqOvRC#DDR8NMRD#CCRO0DHFoOFRVsqR)vnA4_
1cSUz.RH:RVOR5EOFHCH_I8R0E=2RcRMoCC0sNCS
S-V-RHVGRFOsRNRDD4UdU(#,RCODC0VRFRH0s#00NCFRM0CRLHRMosHCo#s0CCS8
RORzE:	RRRHV58N8s8IH0>ERR24.RMoCC0sNCR
RRRRRRORzDR	:bOsFCR##5iBp2R
SRRRRRoLCHSM
RRRRRHRRVBR5pCi'P0CMR8NMRiBpR'=R4R'20MEC
RSRRRRRRRRRNC8so85N8HsI8-0E4FR8IFM0R24.RR<=Ns8_CNo58I8sHE80-84RF0IMF.R42S;
SRRRCRM8H
V;SMSC8sRbF#OC#ORkD
	;SCRRMo8RCsMCNR0Cz	OE;R
RRzRS.:gRRsVFRHHRM8R5CEb0_lMk_DOCD-#RRR428MFI0jFRRMoCC0sNC-
S-VRQR85N8HsI8R0E>.R42CRMC08RFsROCCN0RHIs0CCRMDNLCMRN8kRF00bkRNCMLRDC#CCDOD0RFOoH
RRRRRRRRdSzjRR:H5VRNs88I0H8ERR>4R.2oCCMsCN0
-S-RGVHRsVFRDONDdR4U,U(RD#CCRO0F0VRs0H#NR0CMRF0LMCHoCRso0H#C8sC
RRRRRRRRRRRRRRRR0Fk_5CMH<2R=4R''ERIC5MRNC8so85N8HsI8-0E4FR8IFM0R24.RH=R2DRC#'CRj
';RRRRRRRRRRRRRRRRI_s0CHM52=R<RRW IMECR85N_osC58N8s8IH04E-RI8FMR0F4R.2=2RHR#CDCjR''R;
RRRRRSRRCRM8oCCMsCN0Rjzd;-
S-VRQR85N8HsI8R0E<4=R.M2RFsRIHR0CCLMNDFCRskRF00bkRNCMLRDC#CCDOD0RFOoHRCMC8
C8RRSRRzRSd:4RRRHV58N8s8IH0<ER=.R42CRoMNCs0SC
RRRRRRRRRRRRF_k0CHM52=R<R''4;R
RRRRRRRRRRRRRRsRI0M_C5RH2<W=R R;
RRRRRSRRCRM8oCCMsCN0R4zd;-
S-CRtMNCs00CRE)CRqOvRC#DDR8NMRH0s-N#00
C#RRRRRRRRS.zdRV:RF[sRRRHM58IH0ME_kOl_C#DDR4-R2FR8IFM0RojRCsMCN
0CSNSS0H0sLCk0R_GObbsF#VRFRqA)vj_cgcnXRD:RNDLCRRH#"e1)q"p=R#&RsDPN5[c*+8cRF0IMF*Rc[2+4R"&R,)RWQ_a v m7=&"RR_IslCF8;R
RRRRRRRRRR0RN0LsHkR0C\N3slV_FV0#C\VRFRqA)vj_cgcnXRD:RNDLCRRH#"aA1"RR&HCM0o'CsHolNCH5I820ER"&R7&"RR0HMCsoC'NHloHC5*gcjn&2RR""WRH&RMo0CCHs'lCNo5c[*2RR&"R "&MRH0CCosl'HN5oCo_C0C_M880CbEH55R4+R2j*cgRn,80CbER22&XR""RR&HCM0o'CsHolNC[55+*42c
2;SLSSCMoH
RRRRRRRRRRRR)SAqcv_jXgncRR:)Aqv41n_cR
SRRRRRRRRRbRRFRs0lRNb5R7Q=H>RMC_so*5c[R+d8MFI0cFR*,[2R7q7)>R=RIDF_8N8s454RI8FMR0FjR2, =hR>hR ,1R1)>R=Ra)1,SR
SWSS >R=R0Is_5CMHR2,BRpi=B>RpRi,7dm52>R=R0Fk_#Lkc,5HR[c*+,d2R57m.=2R>kRF0k_L#Hc5,[c*+,.2RS
SSmS75R42=F>RkL0_k5#cH*,c[2+4,mR75Rj2=F>RkL0_k5#cHc,R*2[2;R
RRRRRRRRRRRRRRkRF0C_so*5c[<2R=kRF0k_L#Hc5,[c*2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cco5*4[+2=R<R0Fk_#Lkc,5Hc+*[4I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Coc+*[.<2R=kRF0k_L#Hc5,[c*+R.2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5[c*+Rd2<F=RkL0_k5#cH*,c[2+dRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRCRSMo8RCsMCNR0Cz;d.
RRRRCRSMo8RCsMCNR0Cz;.g
RRRR8CMRMoCC0sNC.RzU
;
SRRRRR--tCCMsCN0RC0ERv)qRDOCDN#RM#8RCODC0FRDoRHOVRFs)Aqv41n_gz
Sd:dRRRHV5FOEH_OCI0H8ERR=go2RCsMCN
0CS-S-RGVHRsVFRDONDdR4U,U(RD#CCRO0F0VRs0H#NR0CMRF0LMCHoCRso0H#C8sC
RSRz	OERH:RVRR5Ns88I0H8ERR>4R42oCCMsCN0
RRRRRRRRDzO	b:RsCFO#5#RB2pi
RSRRRRRLHCoMR
SRRRRRVRHRp5BiP'CCRM0NRM8BRpi=4R''02RE
CMSRRRRRRRRNRR8osC58N8s8IH04E-RI8FMR0F4R42<N=R8C_so85N8HsI8-0E4FR8IFM0R244;S
SRCRRMH8RVS;
S8CMRFbsO#C#RDkO	S;
RMRC8CRoMNCs0zCRO;E	
RRRRdSzcRR:VRFsHMRHRC58b_0EM_klODCD#RR-482RF0IMFRRjoCCMsCN0
-S-RRQV58N8s8IH0>ERR244RCMC8FR0RCOsNR0CI0sHCMRCNCLDR8NMR0FkbRk0CLMND#CRCODC0FRDo
HORRRRRRRRS6zdRH:RVNR58I8sHE80R4>R4o2RCsMCN
0CSR--VRHGVRFsODNDRU4dUR(,#CCDOF0RVsR0HN#00MCRFL0RCoHMRosCHC#0s
C8RRRRRRRRRRRRRRRRF_k0CHM52=R<R''4RCIEMNR58osC58N8s8IH04E-RI8FMR0F4R42=2RHR#CDCjR''R;
RRRRRRRRRRRRRIRRsC0_M25HRR<=WI RERCM5_N8s5CoNs88I0H8ER-48MFI04FR4=2RRRH2CCD#R''j;R
RRRRRRCRSMo8RCsMCNR0Cz;d6
-S-RRQV58N8s8IH0<ER=4R42FRMRHIs0CCRMDNLCsRFR0FkbRk0CLMND#CRCODC0FRDoRHOM8CCCR8
SRRRRdSznRR:H5VRNs88I0H8E=R<R244RMoCC0sNCR
SRRRRRRRRRFRRkC0_M25HRR<=';4'
RRRRRRRRRRRRRRRR0Is_5CMH<2R= RW;R
RRRRRRCRSMo8RCsMCNR0Cz;dn
-S-RMtCC0sNCER0CqR)vCRODRD#NRM80-sH#00NCR#
RRRRRSRRzRd(:FRVsRR[H5MRI0H8Ek_MlC_ODRD#-2R4RI8FMR0FjCRoMNCs0SC
S0SN0LsHkR0CGbO_s#FbRRFVAv)q_c.jURXU:NRDLRCDH"#R1q)epR="&sR#P5NDg+*[gFR8IFM0R[g*+R42&,R"RQW)av _m=7 "RR&Ils_F;8C
RRRRRRRRRRRR0N0skHL0\CR3lsN_VFV#\C0RRFVAv)q_c.jURXU:NRDLRCDH"#RA"1aRH&RMo0CCHs'lCNo58IH0RE2&7R""RR&HCM0o'CsHolNC*5H.Ujc2RR&"RW"&MRH0CCosl'HN5oC[2*gR"&R &"RR0HMCsoC'NHlooC5CC0_M88_CEb05R5H+2R4*c.jU8,RCEb02&2RR""XRH&RMo0CCHs'lCNo5+5[4g2*2S;
SCSLo
HMRRRRRRRRRRRRSqA)vj_.cUUXR):Rq4vAng_1
RSRRRRRRRRRRFRbsl0RN5bR7=QR>MRH_osC5[g*+8(RF0IMF*Rg[R2,q)77RR=>D_FINs885R4j8MFI0jFR2 ,Rh>R=R, hR)11RR=>),1aRS
SS SWRR=>I_s0CHM52B,Rp=iR>pRBi7,Rm25(RR=>F_k0LUk#5UH,*([+27,Rm25nRR=>F_k0LUk#5UH,*n[+2
,RSSSS76m52>R=R0Fk_#LkU,5HU+*[6R2,7cm52>R=R0Fk_#LkU,5HU+*[cR2,7dm52>R=R0Fk_#LkU,5HU+*[dR2,
SSSS57m.=2R>kRF0k_L#HU5,[U*+,.2R57m4=2R>kRF0k_L#HU5,[U*+,42R57mj=2R>kRF0k_L#HU5,[U*2
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRQR7u25jRR=>HsM_Cgo5*U[+27,Rmju52>R=RsbNH_0$LUk#5[H,2
2;RRRRRRRRRRRRRRRRF_k0s5Cog2*[RR<=F_k0LUk#5UH,*R[2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5[g*+R42<F=RkL0_k5#UH*,U[2+4RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_so*5g[2+.RR<=F_k0LUk#5UH,*.[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cgo5*d[+2=R<R0Fk_#LkU,5HU+*[dI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cog+*[c<2R=kRF0k_L#HU5,[U*+Rc2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5[g*+R62<F=RkL0_k5#UH*,U[2+6RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_so*5g[2+nRR<=F_k0LUk#5UH,*n[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cgo5*([+2=R<R0Fk_#LkU,5HU+*[(I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cog+*[U<2R=NRbs$H0_#LkU,5H[I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRS8CMRMoCC0sNCdRz(R;
RRRRS8CMRMoCC0sNCdRzcR;
RCRRMo8RCsMCNR0Cz;dd
R
SR-RR-CRtMNCs00CRE)CRqOvRC#DDR8NMRD#CCRO0DHFoOFRVsqR)vnA4_U14
dSzURR:H5VROHEFOIC_HE80R4=RUo2RCsMCN
0CS-S-RGVHRsVFRDONDdR4U,U(RD#CCRO0F0VRs0H#NR0CMRF0LMCHoCRso0H#C8sC
RSRz	OERH:RVRR5Ns88I0H8ERR>42jRRMoCC0sNCR
RRRRRRORzDR	:bOsFCR##5iBp2R
SRRRRRoLCHSM
RRRRRHRRVBR5pCi'P0CMR8NMRiBpR'=R4R'20MEC
RSRRRRRRRRRNC8so85N8HsI8-0E4FR8IFM0R24jRR<=Ns8_CNo58I8sHE80-84RF0IMFjR42S;
SRRRCRM8H
V;SMSC8sRbF#OC#ORkD
	;SCRRMo8RCsMCNR0Cz	OE;R
RRzRSd:gRRsVFRHHRM8R5CEb0_lMk_DOCD-#RRR428MFI0jFRRMoCC0sNC-
S-VRQR85N8HsI8R0E>jR42CRMC08RFsROCCN0RHIs0CCRMDNLCMRN8kRF00bkRNCMLRDC#CCDOD0RFOoH
RRRRRRRRcSzjRR:H5VRNs88I0H8ERR>4Rj2oCCMsCN0
-S-RGVHRsVFRDONDdR4U,U(RD#CCRO0F0VRs0H#NR0CMRF0LMCHoCRso0H#C8sC
RRRRRRRRRRRRRRRR0Fk_5CMH<2R=4R''ERIC5MRNC8so85N8HsI8-0E4FR8IFM0R24jRH=R2DRC#'CRj
';RRRRRRRRRRRRRRRRI_s0CHM52=R<RRW IMECR85N_osC58N8s8IH04E-RI8FMR0F4Rj2=2RHR#CDCjR''R;
RRRRRSRRCRM8oCCMsCN0Rjzc;-
S-VRQR85N8HsI8R0E<4=RjM2RFsRIHR0CCLMNDFCRskRF00bkRNCMLRDC#CCDOD0RFOoHRCMC8
C8RRSRRzRSc:4RRRHV58N8s8IH0<ER=jR42CRoMNCs0SC
RRRRRRRRRRRRF_k0CHM52=R<R''4;R
RRRRRRRRRRRRRRsRI0M_C5RH2<W=R R;
RRRRRSRRCRM8oCCMsCN0R4zc;-
S-CRtMNCs00CRE)CRqOvRC#DDR8NMRH0s-N#00
C#RRRRRRRRS.zcRV:RF[sRRRHM58IH0ME_kOl_C#DDR4-R2FR8IFM0RojRCsMCN
0CSNSS0H0sLCk0R_GObbsF#VRFRqA)vj_4.4cXnRR:DCNLD#RHR)"1e=qp"RR&#NsPDU54*4[+UFR8IFM0R*4U[2+4R"&R,)RWQ_a v m7=&"RR_IslCF8;R
RRRRRRRRRR0RN0LsHkR0C\N3slV_FV0#C\VRFRqA)vj_4.4cXnRR:DCNLD#RHR1"Aa&"RR0HMCsoC'NHloIC5HE802RR&"R7"&MRH0CCosl'HN5oCHj*4.Rc2&WR""RR&HCM0o'CsHolNC*5[4RU2& R""RR&HCM0o'CsHolNCC5o0M_C8C_8b50E5+HRR*424cj.,CR8b20E2RR&"RX"&MRH0CCosl'HN5oC54[+2U*42S;
SCSLo
HMRRRRRRRRRRRRSqA)vj_4.4cXnRR:)Aqv41n_4RU
RRRRRRRRRRRRRRRRRsbF0NRlb7R5Q>R=R_HMs5Co4[U*+R468MFI04FRU2*[,7Rq7=)R>FRDI8_N8gs5RI8FMR0FjR2, =hR>hR ,1R1)>R=Ra)1,SR
SWSS >R=R0Is_5CMHR2,BRpi=B>RpRi,74m56=2R>kRF0k_L#54nHn,4*4[+6R2,74m5c=2R>kRF0k_L#54nHn,4*4[+cR2,
SSSS57m4Rd2=F>RkL0_kn#454H,n+*[4,d2R57m4R.2=F>RkL0_kn#454H,n+*[4,.2R57m4R42=F>RkL0_kn#454H,n+*[4,42RS
SSmS7524jRR=>F_k0L4k#n,5H4[n*+24j,mR75Rg2=F>RkL0_kn#454H,n+*[gR2,7Um52>R=R0Fk_#Lk4Hn5,*4n[2+U,S
SSmS75R(2=F>RkL0_kn#454H,n+*[(R2,7nm52>R=R0Fk_#Lk4Hn5,*4n[2+n,mR75R62=F>RkL0_kn#454H,n+*[6
2,SRSSR7RRm25cRR=>F_k0L4k#n,5H4[n*+,c2R57md=2R>kRF0k_L#54nHn,4*d[+27,Rm25.RR=>F_k0L4k#n,5H4[n*+,.2
RSSRRRRR7RRm254RR=>F_k0L4k#n,5H4[n*+,42R57mj=2R>kRF0k_L#54nHn,4*,[2RR
RRRRRRRRRRRRRRRRRRRRRRRRRRQR7u>R=R_HMs5Co4[U*+R4(8MFI04FRU+*[4,n2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRu7m5R42=b>RN0sH$k_L#54nH*,.[2+4,mR7u25jRR=>bHNs0L$_kn#45.H,*2[2;R
RRRRRRRRRRRRRRkRF0C_soU54*R[2<F=RkL0_kn#454H,n2*[RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*4[+2=R<R0Fk_#Lk4Hn5,*4n[2+4RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*.[+2=R<R0Fk_#Lk4Hn5,*4n[2+.RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*d[+2=R<R0Fk_#Lk4Hn5,*4n[2+dRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*c[+2=R<R0Fk_#Lk4Hn5,*4n[2+cRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*6[+2=R<R0Fk_#Lk4Hn5,*4n[2+6RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*n[+2=R<R0Fk_#Lk4Hn5,*4n[2+nRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*([+2=R<R0Fk_#Lk4Hn5,*4n[2+(RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*U[+2=R<R0Fk_#Lk4Hn5,*4n[2+URCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*g[+2=R<R0Fk_#Lk4Hn5,*4n[2+gRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*4[+j<2R=kRF0k_L#54nHn,4*4[+jI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co4[U*+244RR<=F_k0L4k#n,5H4[n*+244RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*4[+.<2R=kRF0k_L#54nHn,4*4[+.I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co4[U*+24dRR<=F_k0L4k#n,5H4[n*+24dRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*4[+c<2R=kRF0k_L#54nHn,4*4[+cI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co4[U*+246RR<=F_k0L4k#n,5H4[n*+246RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*4[+n<2R=NRbs$H0_#Lk4Hn5,[.*2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_C4o5U+*[4R(2<b=RN0sH$k_L#54nH*,.[2+4RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRCRSMo8RCsMCNR0Cz;c.
RRRRCRSMo8RCsMCNR0Cz;dg
RRRR8CMRMoCC0sNCdRzU
;
SRRRRR--tCCMsCN0RC0ERv)qRDOCDN#RM#8RCODC0FRDoRHOVRFs)Aqv41n_dSn
zRcd:VRHRE5OFCHO_8IH0=ERR2dnRMoCC0sNCS
S-V-RHVGRFOsRNRDD4UdU(#,RCODC0VRFRH0s#00NCFRM0CRLHRMosHCo#s0CCS8
RORzE:	RRRHV58RN8HsI8R0E>RRg2CRoMNCs0SC
RRRRz	OD:sRbF#OC#BR5p
i2SRSRLHCoMS
SRHRRVBR5pCi'P0CMR8NMRiBpR'=R4R'20MEC
RSSRRRRRsN8CNo58I8sHE80-84RF0IMF2RgRR<=Ns8_CNo58I8sHE80-84RF0IMF2Rg;S
SRCRRMH8RVS;
S8CMRFbsO#C#RDkO	S;
RMRC8CRoMNCs0zCRO;E	
RSRRcRzcRR:VRFsHMRHRC58b_0EM_klODCD#RR-482RF0IMFRRjoCCMsCN0
-S-RRQV58N8s8IH0>ERRRg2M8CCRR0FONsC0ICRsCH0RNCMLRDCNRM8Fbk0kC0RMDNLCCR#D0CORoDFHSO
ScSz6RR:H5VRNs88I0H8ERR>go2RCsMCN
0CSR--VRHGVRFsODNDRU4dUR(,#CCDOF0RVsR0HN#00MCRFL0RCoHMRosCHC#0s
C8SSSSF_k0CHM52=R<R''4RCIEMNR58osC58N8s8IH04E-RI8FMR0Fg=2RRRH2CCD#R''j;S
SSsSI0M_C5RH2<W=R ERIC5MRNs8_CNo58I8sHE80-84RF0IMF2RgRH=R2DRC#'CRj
';SCSSMo8RCsMCNR0Cz;c6
-S-RRQV58N8s8IH0<ER=2RgRRMFI0sHCMRCNCLDRRFsFbk0kC0RMDNLCCR#D0CORoDFHMORCCC88S
SSnzcRH:RVNR58I8sHE80RR<=go2RCsMCN
0CSSSSF_k0CHM52=R<R''4;S
SSsSI0M_C5RH2<W=R S;
SMSC8CRoMNCs0zCRc
n;SR--tCCMsCN0RC0ERv)qRDOCDN#RM08Rs#H-0CN0#S
SS(zcRV:RF[sRRRHM58IH0ME_kOl_C#DDR4-R2FR8IFM0RojRCsMCN
0CSNSS0H0sLCk0R_GObbsF#VRFRqA)v4_6..XdRD:RNDLCRRH#"e1)q"p=R#&RsDPN5*dn[n+dRI8FMR0Fd[n*+R42&,R"RQW)av _m=7 "RR&Ils_F;8C
RRRRRRRRRRRR0N0skHL0\CR3lsN_VFV#\C0RRFVAv)q_.64XRd.:NRDLRCDH"#RA"1aRH&RMo0CCHs'lCNo58IH0RE2&7R""RR&HCM0o'CsHolNC*5H624.R"&RW&"RR0HMCsoC'NHlo[C5*2dnR"&R &"RR0HMCsoC'NHlooC5CC0_M88_CEb05R5H+2R4*.64,CR8b20E2RR&"RX"&MRH0CCosl'HN5oC54[+2n*d2S;
SCSLo
HMSSSSAv)q_.64XRd.:qR)vnA4_n1d
RRRRRRRRRRRRRRRRRRRRRRRRRRRRsbF0NRlb7R5Q>R=R_HMs5Cod[n*+Rd48MFI0dFRn2*[,7Rq7=)R>IDF_8N8sR5U8MFI0jFR2 ,Rh>R=R, hR)11RR=>),1a
SSSSRW =I>RsC0_M25H,pRBi>R=RiBp,mR752d4RR=>F_k0Ldk#.,5Hd[.*+2d4,mR752djRR=>F_k0Ldk#.,5Hd[.*+2dj,S
SSmS752.gRR=>F_k0Ldk#.,5Hd[.*+2.g,mR752.URR=>F_k0Ldk#.,5Hd[.*+2.U,mR752.(RR=>F_k0Ldk#.,5Hd[.*+2.(,S
SSmS752.nRR=>F_k0Ldk#.,5Hd[.*+2.n,mR752.6RR=>F_k0Ldk#.,5Hd[.*+2.6,mR752.cRR=>F_k0Ldk#.,5Hd[.*+2.c,S
SSmS752.dRR=>F_k0Ldk#.,5Hd[.*+2.d,mR752..RR=>F_k0Ldk#.,5Hd[.*+2..,mR752.4RR=>F_k0Ldk#.,5Hd[.*+2.4,S
SSmS752.jRR=>F_k0Ldk#.,5Hd[.*+2.j,mR7524gRR=>F_k0Ldk#.,5Hd[.*+24g,mR7524URR=>F_k0Ldk#.,5Hd[.*+24U,S
SSmS7524(RR=>F_k0Ldk#.,5Hd[.*+24(,mR7524nRR=>F_k0Ldk#.,5Hd[.*+24n,mR75246RR=>F_k0Ldk#.,5Hd[.*+246,S
SSmS7524cRR=>F_k0Ldk#.,5Hd[.*+24c,mR7524dRR=>F_k0Ldk#.,5Hd[.*+24d,mR7524.RR=>F_k0Ldk#.,5Hd[.*+24.,SR
S7SSm4542>R=R0Fk_#LkdH.5,*d.[4+427,Rmj542>R=R0Fk_#LkdH.5,*d.[j+427,Rm25gRR=>F_k0Ldk#.,5Hd[.*+,g2RS
SSmS75RU2=F>RkL0_k.#d5dH,.+*[UR2,7(m52>R=R0Fk_#LkdH.5,*d.[2+(,mR75Rn2=F>RkL0_k.#d5dH,.+*[nR2,
SSSS57m6=2R>kRF0k_L#5d.H.,d*6[+27,Rm25cRR=>F_k0Ldk#.,5Hd[.*+,c2R57md=2R>kRF0k_L#5d.H.,d*d[+2
,RSSSS7.m52>R=R0Fk_#LkdH.5,*d.[2+.,mR75R42=F>RkL0_k.#d5dH,.+*[4R2,7jm52>R=R0Fk_#LkdH.5,*d.[R2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR7RRQ=uR>MRH_osC5*dn[6+dRI8FMR0Fd[n*+2d.,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mud=2R>NRbs$H0_#LkdH.5,[c*+,d2Ru7m5R.2=b>RN0sH$k_L#5d.H*,c[2+.,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mu4=2R>NRbs$H0_#LkdH.5,[c*+,42Ru7m5Rj2=b>RN0sH$k_L#5d.H*,c[;22
RRRRRRRRRRRRRRRRRRRRRRRRFRRks0_Cdo5n2*[RR<=F_k0Ldk#.,5Hd[.*2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRRRRRRRRR0Fk_osC5*dn[2+4RR<=F_k0Ldk#.,5Hd[.*+R42IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[.<2R=kRF0k_L#5d.H.,d*.[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRRRRRRRRR0Fk_osC5*dn[2+dRR<=F_k0Ldk#.,5Hd[.*+Rd2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[c<2R=kRF0k_L#5d.H.,d*c[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRRRRRRRRR0Fk_osC5*dn[2+6RR<=F_k0Ldk#.,5Hd[.*+R62IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[n<2R=kRF0k_L#5d.H.,d*n[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRRRRRRRRR0Fk_osC5*dn[2+(RR<=F_k0Ldk#.,5Hd[.*+R(2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[U<2R=kRF0k_L#5d.H.,d*U[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRRRRRRRRR0Fk_osC5*dn[2+gRR<=F_k0Ldk#.,5Hd[.*+Rg2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[4Rj2<F=RkL0_k.#d5dH,.+*[4Rj2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[4R42<F=RkL0_k.#d5dH,.+*[4R42IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[4R.2<F=RkL0_k.#d5dH,.+*[4R.2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[4Rd2<F=RkL0_k.#d5dH,.+*[4Rd2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[4Rc2<F=RkL0_k.#d5dH,.+*[4Rc2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[4R62<F=RkL0_k.#d5dH,.+*[4R62IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[4Rn2<F=RkL0_k.#d5dH,.+*[4Rn2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[4R(2<F=RkL0_k.#d5dH,.+*[4R(2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[4RU2<F=RkL0_k.#d5dH,.+*[4RU2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[4Rg2<F=RkL0_k.#d5dH,.+*[4Rg2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[.Rj2<F=RkL0_k.#d5dH,.+*[.Rj2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[.R42<F=RkL0_k.#d5dH,.+*[.R42IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[.R.2<F=RkL0_k.#d5dH,.+*[.R.2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[.Rd2<F=RkL0_k.#d5dH,.+*[.Rd2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[.Rc2<F=RkL0_k.#d5dH,.+*[.Rc2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[.R62<F=RkL0_k.#d5dH,.+*[.R62IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[.Rn2<F=RkL0_k.#d5dH,.+*[.Rn2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[.R(2<F=RkL0_k.#d5dH,.+*[.R(2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[.RU2<F=RkL0_k.#d5dH,.+*[.RU2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[.Rg2<F=RkL0_k.#d5dH,.+*[.Rg2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[dRj2<F=RkL0_k.#d5dH,.+*[dRj2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[dR42<F=RkL0_k.#d5dH,.+*[dR42IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[dR.2<b=RN0sH$k_L#5d.H*,c[I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRRRRRRRRRkRF0C_son5d*d[+d<2R=NRbs$H0_#LkdH.5,[c*+R42IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[dRc2<b=RN0sH$k_L#5d.H*,c[2+.RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRRRRRRRRRF_k0s5Cod[n*+2d6RR<=bHNs0L$_k.#d5cH,*d[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''S;
SMSC8CRoMNCs0zCRc
(;SMSC8CRoMNCs0zCRc
c;S8CMRMoCC0sNCcRzd
;
CRM8NEsOHO0C0CksR_MFsOI_E	CO;-

-NRp#H0RlCbDl0CMNF0HM#RHRV8CN0kD
ONsECH0Os0kCCR#D0CO_lsNRRFV)hqv_R)WHV#
k0MOHRFMo_C0C_M880CbEH5#x:CRR0HMCsoCR8;RCEb0RH:RMo0CCRs2skC0sHMRMo0CCHsR#N
PsLHNDlCRH#M_HRxC:MRH0CCos=R:R
j;LHCoMR
Rl_HM#CHxRR:=80CbER;
RRHV5x#HCRR<80CbE02RE
CMRRRRl_HM#CHxRR:=#CHx;R
RCRM8H
V;RCRs0MksRMlH_x#HCC;
Mo8RCC0_M88_CEb0;F
OMN#0MM0RkOl_C#DDRH:RMo0CC:sR=5R55b8C0-ERRR42/.Rd2RR+5855CEb0R4-R2FRl8.Rd2RR/42n2;RRR-y-RRRFV)dqv.1X4RDOCDM#RCCC88OR
F0M#NRM0D0CV_CFPsRR:HCM0oRCs:5=R5C58bR0E+6R42FRl8.Rd2RR/4;n2RRRRRRRRRRRRRRRRRRRRRRRRRR--yVRFRv)q44nX1CRMC88CRsVFRVDC0PRFCIsRF#s8
b0$CkRF0k_L#$_0bHCR#sRNsRN$5lMk_DOCD8#RF0IMF,RjR8IH04E-RI8FMR0FjF2RV0R#8F_Do;HO
o#HMRNDF_k0LRk#:kRF0k_L#$_0bRC;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-7R.RsNsNF$RVFR8k50RHkMb0FR0RH0s-N#002C#
o#HMRNDF_k0C:MRR8#0_oDFHPO_CFO0sk5MlC_ODRD#8MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-MRCNCLD#FRVssR0H0-#N#0C
o#HMRNDF_k0C4M_nRR:#_08DHFoO#;
HNoMDsRI0M_CR#:R0D8_FOoH_OPC05FsM_klODCD#FR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--I0sHCMRCNCLD#FRVsNRCOsERFFIRVqR)vCROD
D##MHoNIDRsC0_Mn_4R#:R0D8_FOoH;H
#oDMNR_HMsRCo:0R#8F_Do_HOP0COFIs5HE80-84RF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-k-R#RC80sFRC#oH0RCs7RQh
o#HMRNDF_k0sRCo:0R#8F_Do_HOP0COFIs5HE80-84RF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-#RkC08RFCRso0H#C7sRm
za#MHoNNDR8C_soRR:#_08DHFoOC_POs0F58N8s8IH04E-RI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RCk#8FR0RosCHC#0s7Rq7#)
HNoMDFRDI8_N8:sRR8#0_oDFHPO_CFO0sR5c8MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--Ns88R0LH#MRHbRk00)FRqOvRC#DDRR5cL#H0RJsCkCHs8N2
0H0sLCk0Rs\3NFl_VCV#0:\RRs#0H;Mo
C
Lo
HM
RRRRR--QNVR8I8sHE80R6<RR#N#HRoM'Rj'0kFRMCk#8HRL0R#
RzRRj:RRRRHV58N8s8IH0=ERRR42oCCMsCN0
RRRRRRRRIDF_8N8s=R<Rj"jjRj"&8RN_osC5;j2
RRRR8CMRMoCC0sNCjRz;R
RR4RzRRR:H5VRNs88I0H8ERR=.o2RCsMCN
0CRRRRRRRRD_FINs88RR<="jjj"RR&Ns8_C4o5RI8FMR0Fj
2;RRRRCRM8oCCMsCN0R;z4
RRRRRz.RH:RVNR58I8sHE80Rd=R2CRoMNCs0RC
RRRRRDRRFNI_8R8s<"=RjRj"&8RN_osC58.RF0IMF2Rj;R
RRMRC8CRoMNCs0zCR.R;
RzRRd:RRRRHV58N8s8IH0=ERRRc2oCCMsCN0
RRRRRRRRIDF_8N8s=R<R''jRN&R8C_soR5d8MFI0jFR2R;
RCRRMo8RCsMCNR0Cz
d;RRRRzRcR:VRHR85N8HsI8R0E>2RcRMoCC0sNCR
RRRRRRFRDI8_N8<sR=8RN_osC58cRF0IMF2Rj;R
RRMRC8CRoMNCs0zCRc
;
RRRR-Q-RV8R5HsM_CRo2sHCo#s0CRh7QRHk#MBoRpRi
RzRR6:RRRRHV5M8H_osC2CRoMNCs0RC
RRRRRbRRsCFO#5#RB,piRh7Q2CRLo
HMRRRRRRRRRRRRH5VRBRpi=4R''MRN8pRBiP'CC2M0RC0EMR
RRRRRRRRRRRRRRMRH_osCRR<=7;Qh
RRRRRRRRRRRR8CMR;HV
RRRRRRRR8CMRFbsO#C#;R
RRMRC8CRoMNCs0zCR6R;
RzRRn:RRRRHV50MFRM8H_osC2CRoMNCs0RC
RRRRRRRRRHRRMC_so=R<Rh7Q;R
RRMRC8CRoMNCs0zCRn
;
RRRR-Q-RV8R5F_k0s2CoRosCHC#0smR7zkaR#oHMRpmBiR
RR(RzRRR:H5VR80Fk_osC2CRoMNCs0RC
RRRRRbRRsCFO#5#RmiBp,kRF0C_soL2RCMoH
RRRRRRRRRRRRRHV5pmBiRR='R4'NRM8miBp'CCPMR020MEC
RRRRRRRRRRRRRRRRz7ma=R<R0Fk_osC;R
RRRRRRRRRRMRC8VRH;R
RRRRRRMRC8sRbF#OC#R;
RRRRRCRRMo8RCsMCNR0Cz
(;RRRRzRUR:VRHRF5M0FR8ks0_CRo2oCCMsCN0
RRRRRRRRRRRRz7ma=R<R0Fk_osC;R
RRMRC8CRoMNCs0zCRU
;
RRRR-Q-RVNR58_8ss2CoRosCHC#0s7Rq7k)R#oHMRiBp
RRRRRzgRH:RVNR58_8ss2CoRMoCC0sNCR
RRRRRRsRbF#OC#BR5pRi,q)772CRLo
HMRRRRRRRRRRRRH5VRBRpi=4R''MRN8pRBiP'CC2M0RC0EMR
RRRRRRRRRRRRRR8RN_osCRR<=q)7758N8s8IH04E-RI8FMR0Fj
2;RRRRRRRRRRRRCRM8H
V;RRRRRRRRCRM8bOsFC;##
RRRR8CMRMoCC0sNCgRz;R
RR4RzjRR:H5VRMRF0Ns88_osC2CRoMNCs0RC
RRRRRRRRRNRR8C_so=R<R7q7)R;
RCRRMo8RCsMCNR0Cz;4j
RRRRRRRRR
RR-R-RMtCC0sNCER0CqR)vCRODRD#NRM8#CCDOD0RFOoH
RRRR4z4RV:RFHsRRRHM5lMk_DOCD-#RRR428MFI0jFRRMoCC0sNCR
RR-R-RRQV58N8s8IH0>ERRR62M8CCRR0FONsC0ICRsCH0RNCMLRDCNRM8Fbk0kC0RMDNLCCR#D0CORoDFHRO
RRRRRzRR4:.RRRHV58N8s8IH0>ERRR62oCCMsCN0
RRRRRRRRRRRRRRRR0Fk_5CMH<2R=4R''ERIC5MRNs8_CNo58I8sHE80-84RF0IMF2R6RH=R2DRC#'CRj
';RRRRRRRRRRRRRRRRI_s0CHM52=R<RRW IMECR85N_osC58N8s8IH04E-RI8FMR0F6=2RRRH2CCD#R''j;R
RRRRRRRRRRMRC8CRoMNCs0zCR4
.;RRRR-Q-RVNR58I8sHE80RR<=6M2RFsRIHR0CCLMNDFCRskRF00bkRNCMLRDC#CCDOD0RFOoHRCMC8
C8RRRRRRRRzR4d:VRHR85N8HsI8R0E<6=R2CRoMNCs0RC
RRRRRRRRRRRRRFRRkC0_M25HRR<=';4'
RRRRRRRRRRRRRRRR0Is_5CMH<2R= RW;R
RRRRRRRRRRMRC8CRoMNCs0zCR4
d;RRRR-t-RCsMCNR0C0REC)RqvODCD#MRN8sR0H0-#N#0C
RRRRRRRRcz4RV:RF[sRRRHM58IH0-ERRR428MFI0jFRRMoCC0sNCR
RRRRRRRRRR0RN0LsHkR0C\N3slV_FV0#C\VRFRqz)vRd.:NRDLRCDH"#R1"1aRH&RMo0CCHs'lCNo58IH0RE2&7R""RR&HCM0o'CsHolNC*5HdR.2&WR""RR&HCM0o'CsHolNC25[R"&R &"RR0HMCsoC'NHlooC5CC0_M88_CEb05R5H+2R4*,d.Rb8C02E2R"&RX&"RR0HMCsoC'NHlo[C5+;42
RRRRRRRRRRRRoLCHRM
RRRRRRRRRzRR)dqv.RR:)dqv.1X4RR
RRRRRRRRRRRRRRFRbsl0RN5bR7>R=R_HMs5Co[R2,q=jR>FRDI8_N8js52q,R4>R=RIDF_8N8s254,.RqRR=>D_FINs885,.2
RRRRRRRRRRRRRRRRRRRRRRRRqRRd>R=RIDF_8N8s25d,cRqRR=>D_FINs885,c2RRW =I>RsC0_M25H,BRWp=iR>pRBim,RRR=>F_k0L5k#H2,[2R;
RRRRRRRRRRRRRFRRks0_C[o52=R<R0Fk_#Lk5[H,2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRCRRMo8RCsMCNR0Cz;4c
RRRRRRRR8CMRMoCC0sNC4Rz4R;RRRRRRRRRRRR
RRRRRR
RR-R-RMtCC0sNCRRN4InRFRs88bCCRv)qRDOCDVRHRbNbssFbHCN0RRRRRRRRRRRRR
RRRRRRzR46:VRHRC5DVF0_PRCs=2R4RMoCC0sNCR
RR-R-RRQV58N8s8IH0>ERRR62M8CCRR0FONsC0ICRsCH0RNCMLRDCNRM8Fbk0kC0RMDNLCCR#D0CORoDFHRO
RRRRRzRR4:nRRRHV58N8s8IH0>ERRR62oCCMsCN0
RRRRRRRRRRRRRRRR0Fk__CM4<nR=4R''ERIC5MR5_N8s5CoNs88I0H8ER-48MFI06FR2RR=M_klODCD#N2RM58RNs8_Cco52RR='2j'2DRC#'CRj
';RRRRRRRRRRRRRRRRI_s0C4M_n=R<RRW IMECRN558C_so85N8HsI8-0E4FR8IFM0RR62=kRMlC_OD2D#R8NMR85N_osC5Rc2=jR''R22CCD#R''j;R
RRRRRRRRRRMRC8CRoMNCs0zCR4
n;RRRR-Q-RVNR58I8sHE80RR<=6M2RFsRIHR0CCLMNDFCRskRF00bkRNCMLRDC#CCDOD0RFOoHRCMC8
C8RRRRRRRRzR4(:VRHR85N8HsI8R0E<6=R2CRoMNCs0RC
RRRRRRRRRRRRRFRRkC0_Mn_4RR<=';4'
RRRRRRRRRRRRRRRR0Is__CM4<nR= RW;R
RRRRRRRRRRMRC8CRoMNCs0zCR4
(;RRRR-t-RCsMCNR0C0REC)RqvODCDR8NMRH0s-N#00RC
RRRRRzRR4:URRsVFRH[RMIR5HE80R4-R2FR8IFM0RojRCsMCN
0CRRRRRRRRRRRRNs00H0LkC3R\s_NlF#VVCR0\FzVR)4qvnRR:DCNLD#RHR1"1a&"RR0HMCsoC'NHloIC5HE802RR&"R7"&MRH0CCosl'HN5oCM_klODCD#.*d2RR&"RW"&MRH0CCosl'HN5oC[&2RR"" RH&RMo0CCHs'lCNo5b8C0RE2&XR""RR&HCM0o'CsHolNC+5[4
2;RRRRRRRRRRRRLHCoMR
RRRRRRRRRR)Rzqnv4R):Rqnv4XR41
RRRRRRRRRRRRRRRRsbF0NRlb7R5RR=>HsM_C[o52q,Rj>R=RIDF_8N8s25j,4RqRR=>D_FINs885,42RRq.=D>RFNI_858s.
2,RRRRRRRRRRRRRRRRRRRRRRRRRdRqRR=>D_FINs885,d2RRW =I>RsC0_Mn_4,BRWp=iR>pRBim,RRR=>F_k0L5k#M_klODCD#2,[2R;
RRRRRRRRRRRRRFRRks0_C[o52=R<R0Fk_#Lk5lMk_DOCD[#,2ERIC5MRF_k0C4M_nRR='24'R#CDCZR''R;
RRRRRRRRRCRRMo8RCsMCNR0Cz;4U
RRRRRRRR8CMRMoCC0sNC4Rz6R;RRRRRRRRR
M
C8sRNO0EHCkO0s#CRCODC0N_sl
;

