--
@ER--B$FbsEHo0OR52gR4g-cRRj.jd$R1MHbDO$H0ROQM
R--fN]C8:CsR#//$DMbH0OH$N/lb..jjDjdNl0/NCbbsN#/0D0/HoL/CFM_s6ONok/lDP03E48yR-f
-


-*-R*************************************************************R**R
---z-RMo#HMRC8v0kDHHbDC-s
-NRas0oCRp:RNH00OmCRsRON6-
-RONsE#DH0RR=DHFoODRLF_O	l0kD
R--4D3RFOoHRN-Rs$sNRDlk0DHbHRCsIEH0RbbHCVLk#HR5MNRO#FCRVHRbbHCDMoHM2-
-
R--.L3RD	FORk-R#oHMROmsNRR6AODF	kRvDb0HDsHCRz5vpUa4X24U

---R-RB$FbsEHo0OR52jR.jRj,.4jjRM1$bODHH,0$ROQM3-
-RDRqDHRso#E0R#sCCCsP8-3
-*R**************************************************************R*R-
-
-*-R*************************************************************R**R
---w-RH0s#u8sFk#O05Rq,Aq,RA-2
--
-R8WH0REq-HRI8R0EFqVRRbHMk-0
-HRW8A0ERI-RHE80RRFVAMRHb
k0-
-R-q-RARR-LIH0NCH#R7qhRRFVNRDDHkMb0-#
--R
-*R**************************************************************R*R-
-
DsHLNRs$HCCC;kR
#HCRC3CC#_08DHFoO4_4nNc3D
D;
LDHs$NsRM#$bVDH$k;
##CR$DMbH3V$Ns00H0LkCN#3D
D;
LDHs$NsROFsN
d;kR#CFNsOds3FOFNOlNb3D
D;
LDHs$NsRM#$bVDH$k;
##CR$DMbH3V$Ns00H0LkCN#3D
D;
0CMHR0$w#Hs0Fus80kO##RH
RRRoCCMs5HO
RRRRIRRHE80qRR:HCM0o;Cs
RRRRIRRHE80ARR:HCM0o
CsR2RR;R
RRsbF0
R5RRRRRRRqRH:RM#RR0D8_FOoH_OPC05FsI0H8E4q-RI8FMR0Fj
2;RRRRRRRARH:RM#RR0D8_FOoH_OPC05FsI0H8E4A-RI8FMR0Fj
2;RRRRRARqRF:Rk#0R0D8_FOoH_OPC05FsI0H8EIA*HE80qR-48MFI0jFR2R
RRRRR-A-RRq*R
RRR2C;
Mw8RH0s#u8sFk#O0;N

sHOE00COkRsCNEsO4VRFRswH#s0uFO8k0H#R#R

RHR#oDMNRNN_k:GRR8#0_oDFHPO_CFO0sH5I8q0E-84RF0IMF2Rj;R
RRo#HMRNDLk_NGRR:#_08DHFoOC_POs0F58IH0-EA4FR8IFM0R;j2
C
Lo
HMRVRRFMsq8Rq:VRFsHHNRMRRj0IFRHE80qR-4oCCMsCN0
RRRRVRRFMsq8RA:VRFsHHLRMRRj0IFRHE80AR-4oCCMsCN0
RRRRRRRRARq58IH0*EAH+NRR2HLRR<=qN5H2hRq75RAH;L2
RRRRCRRMo8RCsMCNR0CVqFsM;8A
RRRCRM8oCCMsCN0RsVFqqM8;M
C8sRNO;E4
-
-R****************************************************************-RR--
-R8N8s5CoqA,R,CR)#-2
--
-RPvFCs#RC#oH0#CsRR0FsDCbNROCbCHbL'kV#-
-R-
-R****************************************************************-RR-D

HNLssH$RC;CCR#
kCCRHC#C30D8_FOoH_n44cD3NDk;
#HCRC3CC#_08DHFoOM_k#MHoCN83D
D;
LDHs$NsRM#$bVDH$k;
##CR$DMbH3V$Ns00H0LkCN#3D
D;
LDHs$NsROFsN
d;kR#CFNsOds3FOFNOlNb3D
D;
0CMHR0$Ns88CHoR#R
RRMoCCOsH5R
RRRRRI0H8ERR:HCM0o;Cs
RRRRsRRCRoRRH:RMo0CC-sR-NRhlFCRVER0CCRDP
CDR2RR;R
RRsbF0
R5RRRRRRRqRRR:H#MR0D8_FOoH_OPC05FsI0H8ER-48MFI0jFR2R;
RRRRRRARRH:RM0R#8F_Do_HOP0COFIs5HE80-84RF0IMF2Rj;R
RRRRR)RC#:kRF00R#8F_Do_HOP0COFIs5HE80-84RF0IMF2Rj
RRR2R;
R0RN0LsHkR0C\N3sMR	\:MRH0CCosR;
R0RN0LsHkR0C\C3slCFP__MFIMNs\RR:HCM0o;Cs
8CMR8N8s;Co
s
NO0EHCkO0sNCRs4OERRFVNs88CHoR#R

RHR#oDMNR#)CkRD0:0R#8F_Do_HOP0COFIs5HE80-84RF0IMF2Rj;L

CMoH
RRR)kC#D<0R=RRq+;RA
RRRVDFsF.Fb:FRVsRRHHjMRRR0FI0H8ER-4oCCMsCN0
RRRRNRR0H0sLCk0Rs\3N\M	RRFVs#CoRD:RNDLCRRH#s;Co
NSS0H0sLCk0Rs\3CPlFCF_M_sINMF\RVCRso:#RRLDNCHDR#;R4
RRRLHCoMR
RRRRRs#Co:HRbbkCLVR
RRRRRb0FsRblN5R
RRRRRRQRRRR=>)kC#DH052R,
RRRRRRRRm>R=R#)C5
H2RRRRR;R2
RRRCRM8oCCMsCN0RsVFDbFF.C;
MN8Rs4OE;-

-*R**************************************************************R*R---
--
-RFVDFQs5M0bk,kRm00bk2-
-
R--****************************************************************R-R-
H
DLssN$CRHCRC;
Ck#RCHCC03#8F_Do_HO4c4n3DND;D

HNLssF$RsdON;#
kCsRFO3NdFNsOObFl3DND;


CHM00V$RDsFFR
H#RoRRCsMCH5OR
RRRRIRRHE80QRhR:MRH0CCos=R:R;dc
RRRRIRRHE80mRza:MRH0CCos=R:R;dc
RRRRMRRkClLsRRR:MRH0CCos=R:R
4;RRRRRMRH8RCGR:RRR0HMCsoCR4:=
RRR2R;
RFRbs50R
RRRRQRRM0bkRRR:RRHM#_08DHFoOC_POs0F58IH0hEQ-84RF0IMF2Rj;R
RRRRRmbk0k:0RR0FkR8#0_oDFHPO_CFO0sH5I8m0Ez4a-RI8FMR0FjR2
R;R2
RRRNs00H0LkC3R\s	NM\RR:HCM0o;Cs
RRRNs00H0LkC3R\sFClPMC_FN_IsRM\:MRH0CCosC;
MV8RDsFF;N

sHOE00COkRsCNEsO4VRFRFVDFHsR#
R
R-RR-CR)o0H#CBsRFFlbM0CM
RRRObFlFMMC08RN8osC
RRRRoRRCsMCH5OR
RRRRRRRRHRI8R0E:MRH0CCosR;
RRRRRRRRsRCoRRR:HCM0oRCs-h-RNRlCF0VREDCRCDPC
RRRR2RR;R
RRRRRb0FsRR5
RRRRRRRRqRRR:MRHR8#0_oDFHPO_CFO0sI5RHE80-84RF0IMF2Rj;R
RRRRRRARRR:RRRRHM#_08DHFoOC_POs0F5HRI8-0E4FR8IFM0R;j2
RRRRRRRRCR)#RR:FRk0#_08DHFoOC_POs0F58IH04E-RI8FMR0FjR2
RRRRR
2;RCRRMO8RFFlbM0CM;R

RHR#oDMNR#)CkRD0:0R#8F_Do_HOP0COFIs5HE80Q4h-RI8FMR0Fj
2;
RRR-V-Rk0MOHRFMONsC0RC#NkRlDb0HDsHCRR0F#VEH0RRNPkNDCCRDVL0R$MRH8RCGL#H0
R
RRMVkOF0HMER#HxV0C5sFHCM8GRR:HCM0o2CsR0sCkRsMHCM0oRCsHR#
RRRRRsPNHDNLC0R#C:bRR0HMCsoC;R
RRoLCHRM
RRRRRC#0b=R:R
4;RRRRRFRVsRRHH4MRRR0FHCM8GR-4DbFF
RRRRRRRR0R#C:bR=0R#C*bRR
.;RRRRRMRC8FRDF
b;RRRRRCRs0MksRC#0bR;
RMRC8ER#HxV0C;sF
R
RRMOF#M0N0ER#HNV08s8CRH:RMo0CC:sR=ER#HxV0C5sFHCM8G
2;RORRF0M#NRM0DoCM0RERR:RRR0HMCsoCRR:=I0H8E/QMMLklC
s;
R--
R--NEsOHO0C0CksRRFVVFDFsRR-FRMCbCHbDCHM80R#N
oC-
-R
oLCH
MRRVRRFFsDF4b_:FRVsRR[H4MRRR0FMLklC.s/RMoCC0sNCR
RRoLCHRM
RRRRRosC#Rq:Ns88CRo
RRRRRMoCCOsHRblNRR5
RRRRRRRRI0H8E>R=RMDCo-0E#VEH08N8C
s,RRRRRRRRRosCR=RR>MRH8
CGRRRRR
R2RRRRRFRbsl0RN
b5RRRRRRRRR=qR>MRQb5k0DoCM05E*.-*[442-RI8FMR0FDoCM0.E**-5[4#2+E0HVNC88s
2,RRRRRRRRR=AR>MRQb5k0DoCM0.E**4[-RI8FMR0FDoCM05E*.-*[4#2+E0HVNC88s
2,RRRRRRRRR#)CRR=>mbk0kD05C0MoE-*[4FR8IFM0RMDCo*0E54[-2E+#HNV08s8C2R
RRRRR2R;
RRRRRsVFDbFF_R.:VRFs	MRHR0jRFER#HNV08s8C-o4RCsMCN
0CRRRRRRRRR0N0skHL0\CR3MsN	F\RVCRso:#RRLDNCHDR#MRH8;CG
SSSNs00H0LkC3R\sFClPMC_FN_IsRM\FsVRCRo#:NRDLRCDH4#R;R
RRRRRLHCoMR
RRRRRR-RR-kRm00bk5MDCo*0E54[-2E+#HNV08s8C-84RF0IMFCRDMEo0*-5[4R22<
=RRRRRRRRRRR--RQRRM0bk5MDCo*0E.[*5-+42#VEH08N8C4s-RI8FMR0FDoCM0.E**-5[4;22
RRRRRRRRCRsoR#:RbbHCVLk
RRRRRRRRFRbsl0RN
b5RRRRRRRRRRRRQ>R=RbQMkD05C0MoE**.54[-22+	,R
RRRRRRRRRRRRm=m>Rkk0b0C5DMEo0*-5[4	2+2R
RRRRRR2RR;R
RRRRRCRM8oCCMsCN0RsVFDbFF_
.;RCRRMo8RCsMCNR0CVDFsF_Fb4
;
RHRRVF_#k:#NRRHV5lMkLRCslRF8.RR=4o2RCsMCN
0CRLRRCMoH
RRRR-RR-sVFDbFF_Rd:VRFsHMRHR04RFCRDMEo0-H#EV80N8RCsoCCMsCN0
RRRRVRRFFsDFdb_:FRVsRRHH4MRRR0FDoCM0oERCsMCN
0CSNSS0H0sLCk0Rs\3N\M	RRFVs#CoRD:RNDLCRRH#HCM8GS;
S0SN0LsHkR0C\C3slCFP__MFIMNs\VRFRosC#RR:DCNLD#RHR
4;RRRRRCRLo
HMRRRRRRRRRosC#R:RbCHbL
kVRRRRRRRRRsbF0NRlbR5
RRRRRRRRRQRRRR=>QkMb0H5I8Q0Eh2-H,R
RRRRRRRRRRRRm=m>Rkk0b0H5I8m0EzHa-2R
RRRRRR2RR;R
RRRRRCRM8oCCMsCN0RsVFDbFF_
d;RRRRR-R-R0mkb5k0I0H8Eamz-H#EV80N8-Cs4FR8IFM0R8IH0zEmaC-DMEo02RR
RRRRRR--R<RR=MRQb5k0I0H8E-Qh#VEH08N8C4s-RI8FMR0FI0H8E-QhDoCM0;E2
RRRCRM8oCCMsCN0R_HV##FkNC;
MN8Rs4OE;-

-*R**************************************************************R*R---
--R
-8RN8aCss5CCR8WH0,EqR8WH02EA
R--
R--****************************************************************R-R-
H
DLssN$CRHCRC;
Ck#RCHCC03#8F_Do_HO4c4n3DND;#
kCCRHC#C30D8_FOoH_HNs0NE3D
D;kR#CHCCC38#0_oDFHkO_Mo#HM3C8N;DD
M
C0$H0R8N8CssaCHCR#R
RRMoCCOsH5R
RRRRRI0H8E:qRR0HMCsoC;R
RRRRRI0H8E:ARR0HMCsoC
RRR2R;
RFRbs50R
RRRRqRRARRRR:RRRRHM#_08DHFoOC_POs0F58IH0*EAI0H8E4q-RI8FMR0Fj
2;RRRRRsRbFO8k0RR:FRk0#_08DHFoOC_POs0F58IH0+EAI0H8E4q-RI8FMR0FjR2
RRRRRR--ARR*qR
RR
2;CRM8NC88sCasCR;

ONsECH0Os0kCsRNORE4FNVR8s8CaCsCR
H#
RRRO#FM00NMRC0EEEHoR#:R0D8_FOoH_OPC05Fs486RF0IMF2RjRR:=Bemh_71a_tpmQeB_ mBa)H5I8q0E-R4,4;n2
R
RRlOFbCFMMV0RDsFF
RRRRoRRCsMCH5OR
RRRRRRRRHRI8Q0Eh:RRR0HMCsoCRR;
RRRRRRRRI0H8EamzRH:RMo0CC;sR
RRRRRRRRkRMlsLCR:RRR0HMCsoCRR;
RRRRRRRRHCM8GRRRRH:RMo0CCRs
RRRRR
2;RRRRRFRbs50R
RRRRRRRRMRQbRk0RH:RM0R#8F_Do_HOP0COFIs5HE80Q4h-RI8FMR0Fj
2;RRRRRRRRR0mkbRk0:kRF00R#8F_Do_HOP0COFIs5HE80m-za4FR8IFM0R
j2RRRRR;R2
RRRCRM8ObFlFMMC0
;
-V-RHRM80RECDNFO0MHFRRFV0RECEEHoCR#0'R4'H"MR0EECH"oE
R
RRMVkOF0HMCR8bW0EHE80R0sCkRsMHCM0oRCsHR#
RCRLo
HMRRRRRFRVsRRHH4MR6FR8IFM0RDjRF
FbRRRRRRRRRRHV5C0EEEHo5RH2=4R''02RE
CMRRRRRRRRRRRRR0sCkRsMH;+4
RRRRRRRRMRC8VRH;R
RRRRRCRM8DbFF;R
RRRRRskC0sjMR;R
RR8CMRb8C0HEW8;0E
R
RRMOF#M0N0CR8bR0ERH:RMo0CC:sR=CR8bW0EHE80;R
RRMOF#M0N0HRI8R0E:MRH0CCos=R:R8IH0+EAI0H8E4q+;R
RRb0$CHRDlH#R#sRNsRN$5b8C04E+RI8FMR0FjF2RVMRH0CCosR;

R--V8HMRC0ERJsCkCHs8kRMlsLC#0R5EMC_kClLsH#RMMRNRsNsNF$RVMRH0CCos
#2
RRRVOkM0MHFRDONOlhkL#CsR0sCkRsMD#HlR
H#RRRRRNRPsLHND0CREMC_kClLs:#RRlDH#R;
RCRLo
HMRRRRRER0Ck_MlsLC#25jRR:=I0H8E
q;RRRRRFRVsRRHH4MRRR0F80CbER+4DbFF
RRRRRRRRER0Ck_MlsLC#25HRR:=0_ECMLklC5s#H2-4/+.RRE50Ck_MlsLC#-5H4l2RF.8R2R;
RRRRR8CMRFDFbR;
RRRRR0sCkRsM0_ECMLklC;s#
RRRR8CMRDONOlhkL#Cs;

RRORRF0M#NRM0MLklCRs#:HRDl:#R=NRODkOhlsLC#R;

R--OONDk0DNCER0CH_Dl
#
RVRRk0MOHRFMOONDpRHlskC0sDMRHRl#HR#
RRRRRsPNHDNLCER0CH_Dl:#RRlDH#R;
RRRRRsPNHDNLCkRMlRLRR:RRR0HMCsoC;R
RRoLCHRM
RRRRRC0E_lDH#25jRR:=jR;
RRRRRlMkL=R:R8IH0;Eq
RRRRVRRFHsRRRHM4FR0Rb8C04E+RFDFbR
RRRRRR0RREDC_H5l#H:2R=ER0CH_DlH#5-R42+kRMlIL*HE80;R
RRRRRRMRRkRlL:M=Rk/lL.RR+5lMkLFRl82R.;R
RRRRRCRM8DbFF;R
RRRRRskC0s0MREDC_H;l#
RRRCRM8OONDp;Hl
RR
RFROMN#0MP0RCHODlRR:D#HlRR:=OONDp;Hl
RRR#MHoNRDRL0HosRCC:0R#8F_Do_HOP0COFPs5CHODlC58b+0E442-RI8FMR0Fj
2;
R--ONsC00CRENCRsHOE00COkRsCF0VRENCR8s8CRC0sCL

CMoHRR
RRsVFNqM8:FRVsNRHRRHMjFR0R8IH0-Eq4CRoMNCs0RC
RRRRRoLH0CsC5N5H+*42I0H8ER-48MFI0HFRNH*I820ERR<=RhBmea_17m_pt_QBea Bmj)5,HRI8q0E-+HN4R2
RRRRRRRR&ARq58IH0*EA5+HN442-RI8FMR0FI0H8EHA*NR2
RRRRRRRR&mRBh1e_ap7_mBtQ_Be a5m)jH,RN
2;RCRRMo8RCsMCNR0CVNFsM;8q
R
RRsVFDbFF.F:VsRR[H4MRRR0F80CbECRoMNCs0RC
R4Rl:VRRDsFF
RRRRoRRCsMCHlORN5bR
RRRRRRRRHRI8Q0Eh=RR>CRPOlDH5R[2-CRPOlDH54[-2R,
RRRRRRRRI0H8EamzRR=>PDCOH[l5+R42-CRPOlDH5,[2
RRRRRRRRkRMlsLCR=RR>kRMlsLC#-5[4
2,RRRRRRRRR8HMCRGRR>R=RR[
RRRRRRRR2R
RRRRRb0FsRblNRR5
RRRRRRRRQkMb0RRRRR=>L0Hos5CCPDCOH[l52R-48MFI0PFRCHODl-5[4,22
RRRRRRRRkRm00bkR=RR>HRLoC0sCC5POlDH54[+2R-48MFI0PFRCHODl25[2R
RRRRR2R;
RMRC8oRRCsMCNR0CVDFsF.Fb;R

RsRbFO8k0=R<RoLH0CsC5OPCD5Hl80CbE2+4-8.RF0IMFCRPOlDH5b8C02E2;
R
CRM8NEsO4
;
-*-R*************************************************************
**-a-REkCRMo#HMRC8l0kDH$bDRCk##zRvp(a4G
4(-*-R*************************************************************
**
LDHs$NsR Q  k;
#HCRC3CC#_08DHFoO4_4nNc3D
D;kR#CHCCC38#0_oDFHNO_sEH03DND;#
kCCRHC#C30D8_FOoH_o#HM3C8N;DD
M
C0$H0RpvzaX4(4H(R#

SRbRRFRs05R
RRRRRqRR:HRMR#_08DHFoOC_POs0F5R4n8MFI0jFR2R;
RRRRR:ARRRHMR8#0_oDFHPO_CFO0sn54RI8FMR0Fj
2;RRRRRRRu:kRF00R#8F_Do_HOP0COFds5dFR8IFM0R
j2S;S2
R
RR0N0skHL0\CR30HMCNsMDM_H#M0N00HNCR8\:MRH0CCosC;
Mv8Rz4pa((X4;-

-$R#MC0E#RH#0MsN#0DNCV_FV-
-RLDHs$NsRl#HblsH;-
-RCk#Rl#HblsH3NebOo	NCD3ND-;
-$R#MC0E#RH#0MsN#0DNCM_F
s
NO0EHCkO0s#CR0Osk0VRFRpvzaX4(4H(R#R

RFROlMbFCRM0vazp44UXUv_ 
RRRRbRRFRs05S
Sq,4(Rnq4,4Rq6q,R4Rc,q,4dR.q4,4Rq4q,R4Rj,qRgRRRRRR:RRRRHM#_08DHFoO
R;SUSq,(Rq,nRq,6Rq,cRq,dRq,.Rq,4Rq,jRqSSSSR:RRRRHM#_08DHFoO
R;S4SA(A,R4Rn,A,46RcA4,4RAdA,R4R.,A,44RjA4,gRARRRRRRRRRH:RM0R#8F_DoRHO;S
SARU,AR(,ARn,AR6,ARc,ARd,AR.,AR4,ASjSSRSRRH:RM0R#8F_DoRHO;S

RRRRu,d6Rcud,dRudu,RdR.,u,d4Rjud,.Rugu,R.RU,uR.(RRRRR:RRR0FkR8#0_oDFH;OR
uSS.Rn,u,.6Rcu.,.Rudu,R.R.,u,.4Rju.,4Rugu,R4SUSR:RRR0FkR8#0_oDFH;OR
uSS4R(,u,4nR6u4,4Rucu,R4Rd,u,4.R4u4,4Ruju,RgRRRRRRRRRR:FRk0#_08DHFoO
R;SUSu,(Ru,nRu,6Ru,cRu,dRu,.Ru,4Ru,jRuSSSSR:RRR0FkR8#0_oDFH
ORS;S2
MSC8FROlMbFC;M0
R
RR0N0skHL0#CR$LM_D	NO_GLFRL:RFCFDN
M;RNRR0H0sLCk0RM#$_NLDOL	_FFGRVzRvpUa4X_4U :vRRlOFbCFMMH0R#)Raz
 ;
HS#oDMNRhqQR#:R0D8_FOoH_OPC0RFs5R4(8MFI0jFR2S;
#MHoNADRQ:hRR8#0_oDFHPO_CFO0s4R5(FR8IFM0R;j2
#
SHNoMD)Rum:7RR8#0_oDFHPO_CFO0sdR56FR8IFM0R;j2
N
S0H0sLCk0RH\3Ms0CM_NDH0M#NHM0N80C\VRFRDlk0RR:DCNLD#RHR
4;LHCoMR

RQRqh=R<R""jRq&R;-SR-kRb0RRNxFCsRRHMVMsF0R
RRhAQRR<="Rj"&;RA
l
SkRD0:zRvpUa4X_4U Rv
RRRRRsbF0NRlb
R5RRRRRRRRRqRR4=(R>QRqh(542R,
RRRRRRRRqR4n=q>RQ4h5n
2,RRRRRRRRR6q4RR=>q5Qh4,62
RRRRRRRR4Rqc>R=RhqQ524c,R
RRRRRRqRR4=dR>QRqhd542R,
RRRRRRRRqR4.=q>RQ4h5.
2,RRRRRRRRR4q4RR=>q5Qh4,42
RRRRRRRR4Rqj>R=RhqQ524j,R
RRRRRRqRRg>R=RhqQ5,g2
RRRRRRRRURqRR=>q5QhU
2,RRRRRRRRRRq(=q>RQ(h52R,
RRRRRRRRq=nR>QRqh25n,R
RRRRRRqRR6>R=RhqQ5,62
RRRRRRRRcRqRR=>q5Qhc
2,RRRRRRRRRRqd=q>RQdh52R,
RRRRRRRRq=.R>QRqh25.,R
RRRRRRqRR4>R=RhqQ5,42
RRRRRRRRjRqRR=>q5Qhj
2,RRRRRRRRR(A4RR=>A5Qh4,(2
RRRRRRRR4RAn>R=RhAQ524n,R
RRRRRRARR4=6R>QRAh6542R,
RRRRRRRRAR4c=A>RQ4h5c
2,RRRRRRRRRdA4RR=>A5Qh4,d2
RRRRRRRR4RA.>R=RhAQ524.,R
RRRRRRARR4=4R>QRAh4542R,
RRRRRRRRAR4j=A>RQ4h5j
2,RRRRRRRRRRAg=A>RQgh52R,
RRRRRRRRA=UR>QRAh25U,R
RRRRRRARR(>R=RhAQ5,(2
RRRRRRRRnRARR=>A5Qhn
2,RRRRRRRRRRA6=A>RQ6h52R,
RRRRRRRRA=cR>QRAh25c,R
RRRRRRARRd>R=RhAQ5,d2
RRRRRRRR.RARR=>A5Qh.
2,RRRRRRRRRRA4=A>RQ4h52R,
RRRRRRRRA=jR>QRAh25j,R
RRRRRRuRRd=6R>)Rumd756
2,RRRRRRRRRcudRR=>u7)m52dc,R
RRRRRRuRRd=dR>)Rumd75d
2,RRRRRRRRR.udRR=>u7)m52d.,R
RRRRRRuRRd=4R>)Rumd754
2,RRRRRRRRRjudRR=>u7)m52dj,R
RRRRRRuRR.=gR>)Rum.75g
2,RRRRRRRRRUu.RR=>u7)m52.U,R
RRRRRRuRR.=(R>)Rum.75(
2,RRRRRRRRRnu.RR=>u7)m52.n,R
RRRRRRuRR.=6R>)Rum.756
2,RRRRRRRRRcu.RR=>u7)m52.c,R
RRRRRRuRR.=dR>)Rum.75d
2,RRRRRRRRR.u.RR=>u7)m52..,R
RRRRRRuRR.=4R>)Rum.754
2,RRRRRRRRRju.RR=>u7)m52.j,R
RRRRRRuRR4=gR>)Rum475g
2,RRRRRRRRRUu4RR=>u7)m524U,R
RRRRRRuRR4=(R>)Rum475(
2,RRRRRRRRRnu4RR=>u7)m524n,R
RRRRRRuRR4=6R>)Rum4756
2,RRRRRRRRRcu4RR=>u7)m524c,R
RRRRRRuRR4=dR>)Rum475d
2,RRRRRRRRR.u4RR=>u7)m524.,R
RRRRRRuRR4=4R>)Rum4754
2,RRRRRRRRRju4RR=>u7)m524j,R
RRRRRRuRRg>R=Rmu)725g,R
RRRRRRuRRU>R=Rmu)725U,R
RRRRRRuRR(>R=Rmu)725(,R
RRRRRRuRRn>R=Rmu)725n,R
RRRRRRuRR6>R=Rmu)7256,R
RRRRRRuRRc>R=Rmu)725c,R
RRRRRRuRRd>R=Rmu)725d,R
RRRRRRuRR.>R=Rmu)725.,R
RRRRRRuRR4>R=Rmu)7254,R
RRRRRRuRRj>R=Rmu)725j
2SS;S
S
RRRu=R<Rmu)7d5dRI8FMR0FjS2;RR--0CN	RDFM$cRdR0LH#C

M#8R0Osk0
;
-*-R*************************************************************R**R
---e-R.mApBqi5,,RARmu)7-2
--
-RHNI8R0E-HRI8R0EFqVRRbHMk-0
-IRLHE80RI-RHE80RRFVAMRHb
k0-
-R-u-R)Rm7-ERaCkRVDbDRskF8O50RN8IH0+ERRHLI8R0EICH82sRVFLlRD	FORDlk0DHbH#Cs3-R
--R
-*R**************************************************************R*R-
-
DsHLNRs$HCCC;#
kCCRHC#C30D8_FOoH_n44cD3NDk;
#HCRC3CC#_08DHFoOs_NH30EN;DD
Ck#RCHCC03#8F_Do_HOkHM#o8MC3DND;D

HNLssF$RsdON;#
kCsRFO3NdFNsOObFl3DND;C

M00H$.ReABpmi#RH
CSoMHCsO
R5SISNHE80RH:RMo0CC
s;SISLHE80RH:RMo0CC
s;SCSMCb8_HDbCHRMC:MRH0CCos2
S;b
SFRs05S
SqRRRRH:RM#RR0D8_FOoH_OPC05FsN8IH04E-RI8FMR0Fj
2;SRSAR:RRRRHMR8#0_oDFHPO_CFO0sI5LHE80-84RF0IMF2Rj;S
Su7)mRF:Rk#0R0D8_FOoH_OPC05FsN8IH0LE+I0H8ER-48MFI0jFR22
S;N
S0H0sLCk0Rs\3N\M	RH:RMo0CC
s;S0N0skHL0\CR3oLCH0M_s\CCRH:RMo0CC
s;S0N0skHL0\CR3lsCF_PCMIF_N\sMRH:RMo0CC
s;CRM8ep.Am;Bi
s
NO0EHCkO0sLCRD	FO#VRFRAe.pimBR
H#
-S-RlqRNlGHkVlRk0MOHRFMM8CCCI8RERCMN8IH0HER#FRM0JRCkRND0LFRI0H8E-
S-kRbs#bFCV:RHRM80REC#NJksNCRs$sNR8IH0VERsRFl0RECHkMb0kRL#HR#x
C#RVRRk0MOHRFMlN$lGPR5NCDkNP,RNCDkLRR:HCM0o2Cs
sSSCs0kMMRH0CCos#RH
CSLoRHMRR--lN$lGS
SHPVRNCDkNRR>PkNDC0LRE
CMSsSSCs0kMNRPDNkC;S
SCCD#
SSSskC0sPMRNCDkLS;
S8CMR;HV
MSC8$Rll;NG
R
RRlOFbCFMMv0Rz4pa((X4
RRRRbRRFRs05R
RRRRRRqRRRH:RM#RR0D8_FOoH_OPC0RFs5R4n8MFI0jFR2R;
RRRRRRRRARR:HRMR#_08DHFoOC_POs0FRn54RI8FMR0Fj
2;RRRRRRRRR:uRR0FkR8#0_oDFHPO_CFO0sdR5dFR8IFM0R
j2S;S2
RRRCRM8ObFlFMMC0
;
RORRF0M#NRM0WRzvR:RRR0HMCsoCRR:=4
(;
RRRO#FM00NMR)Z mR4(:0R#8F_Do_HOP0COF:sR=jR"jjjjjjjjjjjjjjjj"
;
SMOF#M0N0HRI8RNRRH:RMo0CC:sR=5R5N8IH0WE+z4v-2z/Wv
2;RORRF0M#NRM0ILH8R:RRR0HMCsoCRR:=5I5LHE80+vWz-/42W2zv;R
RRMOF#M0N0bRIsR8RRH:RMo0CC:sR=HRI8+NRR8IHLS;
O#FM00NMRsINsRRR:MRH0CCos=R:R8IHNRR*ILH8;R
RRMOF#M0N0lRINRGRRH:RMo0CC:sR=$Rll5NGINH8,HRI8;L2
-
S-ERaCMRHb#k0RCNsRD#bHH0RMR0F4L(-HO0RE	kM#R
RRb0$C0Rq$RbCHN#Rs$sNRR5j0IFRH-8N4F2RV0R#8F_Do_HOP0COFRs5RvWz-84RF0IMF2Rj;R
RRb0$C0RA$RbCHN#Rs$sNRR5j0IFRH-8L4F2RV0R#8F_Do_HOP0COFRs5RvWz-84RF0IMF2Rj;S

-0-RECCRDCClMR0#F0VREuCRNHs0N1DRk)lRFRI#NRsC4L(-HR0#ICH8
$S0b1CR0C$bRRH#NNss$jR5RR0FI8bs-R42F#VR0D8_FOoH_OPC05FsRzRWvR-48MFI0jFR2
;
SR--0RECb0NsHRNDb8sFk#O0RCNsR-dcL#H0R8IHC.R5*vWz20
S$RbCub0$C#RHRsNsN5$RjFR0RsINs2-4RRFV#_08DHFoOC_POs0F5W.*z4v-RI8FMR0Fj
2;
-S-RCaERbHMkR0#HNMRR8IHNsRNsRN$F4VRUH-L0EROk#M	
HS#oDMNRsqNsRN$R:RRR$q0b
C;So#HMRNDAsNsNR$RRRR:Ab0$C
;
SR--0RECu0NsHRNDu8sFkRO0NNss$#RNRINRNRssNNss$VRFR-dnLRH0OMEk	R#
RHR#oDMNRkuLVRRRR:RRR$u0b
C;R#RRHNoMDsRuFs8qsRN$:0Ru$;bC
LS
CMoHR-R-RFLDOl	_k
D0
-S-RCaE#0CRIbFRsCFO###CRNOEMRoC0RECPHNsNCLDR8IH0HERM0bk#MRH0VFRH8GCR8IH0HERM0bk#S3
-a-REICRHE80RRFV0RECHkMb0N#RsHCRMzRWvsRoF#kbRsVFR0LFER3
RCRs#CHx_RN:bOsFCR##5Rq,qsNsN
$2SoLCHRMR-b-RsCFO#s#RCx#HC
_NSNSqs$sN58IHN2-4RR<= 5XaqI5NHE80-84RF0IMFzRWvI*5H-8N4,22RvWz2S;
SsVFRGH8RRHMjFR0R8IHNR-.DbFF
SSSqsNsNH$58RG2<q=R5vWz*85HG2+4-84RF0IMFzRWv8*HG
2;RRRRRMRC8FRDF
b;S8CMRFbsO#C#R#sCH_xCN
;
RsRRCx#HC:_LRFbsO#C#R,5ARsANs2N$
RRRLHCoM-RR-sRbF#OC#CRs#CHx_SL
SsANs5N$ILH8-R42< =RXAa55HLI8-0E4FR8IFM0RvWz*H5I84L-2R2,W2zv;R
RRRRRVRFsHR8GHjMRRR0FILH8-D.RF
FbSASSNNss$85HG<2R=5RAW*zv5GH8+-424FR8IFM0RvWz*GH82S;
S8CMRFDFbR;R-H-R8RG
RMRC8sRbF#OC#CRs#CHx_
L;
-S-RMoCC0sNCER0CNRusN0HDsRuFO8k0sRNsRN$Ll$RkHD0bHD$M0oRE4CRUH-L0EROk#M	R
FVSR--0RECHkMb00#RFFRVsdlRnH-L0NRusN0HDsRuFO8k0R#3RR

RCRoMDlk0RN:VRFsNHGRMRRj0IFRH-8N4CRoMNCs0SC
SMoCl0kDLV:RFLsRGMRHR0jRFHRI84L-RMoCC0sNCS
SSDlk0:GRRpvzaX4(4S(
SbSSFRs0lRNb5S
SSqSSRR=>qsNsNN$5G
2,SSSSS=AR>NRAs$sN52LG,S
SSuSSRR=>uVLk5G5N*8IHLL2+GS2
SSSS2S;
SVSH_bbHNR4:H5VRM8CC_bbHCMDHCRR=4o2RCsMCN
0CSSSSLbkVbRH:VRFsHMRHR0jRF*R.W-zv4CRoMNCs0SC
SSSSNs00H0LkC3R\s	NM\VRFRosC#RR:DCNLD#RHR
4;SSSSS0N0skHL0\CR3oLCH0M_s\CCRRFVs#CoRD:RNDLCRRH#4S;
SSSSNs00H0LkC3R\sFClPMC_FN_IsRM\FsVRCRo#:NRDLRCDH4#R;S
SSCSLoRHM
SSSSCSsoR#:RbbHCVLk
SSSSbSSFRs0l5Nb
SSSSSSSQ>R=RkuLVN55GH*I8+L2L5G2H
2,SSSSSmSSRR=>u8sFqNss$N55GH*I8+L2L5G2HS2
SSSSS
2;SSSSCRM8oCCMsCN0RVLkb;bH
SSSCRM8oCCMsCN0R_HVbNHb4S;
SVSH_bbHNRj:H5VRM8CC_bbHCMDHCRR=jo2RCsMCN
0CSSSSu8sFqNss$N55GH*I8+L2LRG2<u=RL5kV5*NGILH82G+L2S;
SMSC8CRoMNCs0HCRVH_bb;Nj
CSSMo8RCsMCNR0ColCMkLD0;C
SMo8RCsMCNR0ColCMkND0;S

-a-RNR	C0RECu0NsHRNDu8sFkRO0NNss$MRN8kRLHRD80RECNC88ssR0CRC3RsqRkHMMM#oRkSl
-H-R#MRHHD0NH8xC,ER0CFMR0sECRIsF#VRFRC0ERsbN0DHNRFbs80kORCNsR8N8C
83SR--wRFsClGNb,DCRRHVq#RHR-6UL#H0R8IHCMRN8RRAH.#RcH-L0I#RH,8CRC0EMRRqV#H0RRHMc-
S-(R4-0LHRkOEMR	#NRM8AHRV0H#RMRR.4L(-HO0RE	kM#R3RaRECNNss$HRIDHDRMkOD8cCR*
.=SR--UkRlDb0HDsHC#FRVsMlHoRRUdLn-Hu0RNHs0NuDRskF8O30#RERaCkRVDbDRskF8OI0RHRDDL
CRSR--c=+.n(R4-0LHRkOEMR	#ICH83wRRF0sRERH#ClGNbRDC0REC)1kMkHlR#MRHHN0HDCHx8FR0:-
S-RRRR#j',RRRRRRRj,'#RRRRRuRRu,544H2E,uRu544,2,DFR5uuj2,jERH,uju5,Dj2F-
S-ERaCFMR0sECRIsF#sRNCFRVs8lCR#LNCF8RMER0CHRI8R0EFqVRRRHM4L(-HO0RE	kM#MRN8-
S-ER0CHRI8R0EFAVRRRHM4L(-HO0RE	kM#R3RwRFs0RECClGNb:DC
-S-RCaER''qRFDFb4R5RR0FdS2
-R-RR'Rj#R,RRRRRR5uu.2,4ERH,u.u5,D42Fu,Ru,54jH2E,uRu5j4,2,DFR#j'
-S-RRRRudu5,E42Hu,Ru,5d4F2D,uRu5j.,2,EHR5uu.2,jDRF,j,'#RRRRRjRR'S#
-R-RR'Rj#R,RRRRRR5uud2,jERH,udu5,Dj2Fj,R'R#,RRRRR'Rj#R,RRRRRR#j'
-S-RCaER''ARFDFb4R5RR0F4S2
-R-RR'Rj#R,RRRRRR#j',RRRRRRRj,'#RRRRRuRRu,5j4H2E,uRu54j,2,DFR#j'
R
RR8N8b8sF:sRbF#OC#uR5sqF8s$sN2S
SPHNsNCLDRM)k1RklR:RRR8#0_oDFHPO_CFO0sb5IsW8*z4v-RI8FMR0Fj:2R=FR50sEC#>R=R''j2R;
RRRRRsPNHDNLCkR1lI)FeRCO:0R#8F_Do_HOP0COFIs5b*s8W-zv4FR8IFM0R;j2
RRRRPRRNNsHLRDC1)klFRIRRRR:1b0$CR;
RRRRRsPNHDNLCHRN8RGRRRRR:MRH0CCosR;
RRRRRsPNHDNLCHRL8RGRRRRR:MRH0CCosR;
RRRRRsPNHDNLCRR[RRRRRRRR:MRH0CCosR;
RRRRRsPNHDNLCRR	RRRRRRRR:MRH0CCosS;
LHCoM-RR-sRbF#OC#8RN8Fbs8S
S-Q-RMHH0NxDHCER0CkRsMMMHokR#l)R5kkM1lR2
RRRRRsVFRRNGHjMRRR0FIGlN-D4RF
FbSLSSHR8G:N=RGS;
SRS[R:RR=*R.N
G;S	SSRRRR:[=RR4+R;S
SSRHVN>GRR8IHNR-4FLsRHR8G>HRI84L-RC0EMS
SSVSHR<[RRsIb8ER0CRMRS-SR-CRxsCFRGM0C8S
SS1SSkFl)I25[RR:=Zm )4
(;SSSSCRM8H
V;SSSSH	VRRI<RbRs80MECRSRSRR--xFCsR0CGC
M8SSSSSl1k)5FI	:2R= RZ)(m4;S
SSMSC8VRH;S
SS#CDCS
SSkS1lI)F5R[2:u=RsqF8s$sN5*NGILH8+8LHGR25RvWz-84RF0IMFRRRj
2;RRRRRRRRRRRRH	VRRI<RbRs80MEC
SSSSkS1lI)F5R	2:u=RsqF8s$sN5*NGILH8+8LHG.25*vWz-84RF0IMFzRWv
2;SSSSCRM8H
V;SCSSMH8RVS;
S-S-RMOFP0CsRC0ERsNsNF$RVEROk#M	R0HMFMRNRsNsNF$RVHRL0S#
SFSVsLRHGMRHR0jRFbRIs48-RFDFbS
SSFSVsGRDRRHMjFR0RvWz-D4RF
FbSSSSSM)k15klH*LGW+zvDRG2:1=RkFl)IL5HGD25G
2;SSSSCRM8DbFF;-RR-GRD
SSSCRM8DbFF;-RR-LRHGS
SCRM8DbFF;-RR-GRN
-SS-FRpFFbRMER0CRRqHCM8GS
SVRFsHR8GH4MRRR0FINH8-D4RF
FbRRRRRRRRRsVFRRNGHjMRRR0FIGlN-D4RF
FbSSSSLGH8RR:=N-GRRGH8;S
SSRS[R:RR=GRNRL+RH;8G
SSSSR	RR=R:R+[RR
4;SSSSHNVRGRR>INH8-F4RsHRL8>GRR8IHLR-40MEC
RRRRRRRRRRRRRRRH[VRRI<RbRs80MECRSRSRR--xFCsR0CGC
M8SSSSSkS1lI)F5R[2:Z=R 4)m(S;
SSSSCRM8H
V;SSSSSRHV	RR<I8bsRC0EMSRRS-R-RsxCFGRC08CM
SSSS1SSkFl)I25	RR:=Zm )4
(;SSSSS8CMR;HV
SSSS#CDHLVRHR8G<RRj0MEC
SSSSVSHR<[RR0jRE
CMSSSSSRS[:[=RR.+R*NIlGR;
RRRRRRRRRRRRRMRC8VRH;R
RRRRRRRRRRRRRRRHV	RR<jER0CSM
SSSSS:	R=RR	+*R.IGlN;S
SSCSSMH8RVS;
SSSSH[VRRN<RGER0CSM
SSSSSl1k)5FI[:2R= RZ)(m4;S
SSCSSDV#HR<[RRsIb8ER0CSM
SSSSSl1k)5FI[:2R= RZ)(m4;-RR-CRxsCFRGM0C8S
SSCSSMH8RVS;
SSSS-F-R0sECICH#,ER0CMRH8RCGHM#RFH0RMER0CkR1lI)F,FR8R0MFEoHM
SSSSVSHR<	R=GRNRC0EMS
SSSSS1)klF	I52=R:R)Z m;4(
RRRRRRRRRRRRRRRCHD#VRR	<bRIs08RE
CMSSSSSkS1lI)F5R	2:Z=R 4)m(R;R-x-RCRsFCCG0MS8
SSSS-F-R0sECICH#,ER0CMRH8RCGHM#RFH0RMER0CkR1lI)F,FR8R0MFEoHM
SSSSMSC8VRH;S
SSDSC#SC
SSSS1)klF[I52=R:RFus8sqsNN$5GH*I8LL+H28G5WRRz4v-RI8FMR0FR2Rj;R
RRRRRRRRRRRRRRRHV	RR<I8bsRC0EMS
SSSSS1)klF	I52=R:RFus8sqsNN$5GH*I8LL+H28G5W.*z4v-RI8FMR0FW2zv;S
SSCSSMH8RVS;
SCSSMH8RVS;
SMSC8FRDFRb;RR--NSG
S-S-RMOFP0CsRC0ERsNsNF$RVEROk#M	R0HMFMRNRsNsNF$RVHRL0R#
RRRRRRRRVRFsHRLGHjMRRR0FI8bs-D4RF
FbSSSSVRFsDHGRMRRj0WFRz4v-RFDFbS
SS1SSkFl)IOeC5GHL*vWz+2DGRR:=1)klFHI5L5G2D;G2
SSSS8CMRFDFbR;R-D-RGS
SS8CMRFDFbR;R-H-RLSG
S-S-R8q8RC0ERIsFR#[k0sROCCN08FR0RC0ERMskMoHMRl#k
RRRRRRRRkR)Ml1kRR:=)1kMk+lRRl1k)eFIC
O;SMSC8FRDFRb;RR--H
8GS-S-RFpFbMRFRC0ERHARMG8C
VSSFHsRxHGRMRR40IFRH-8L4FRDFRb
RRRRRRRRVRFsLHGRMRRj0IFRl-NG4FRDFSb
SNSSHR8G:L=RGRR-H;xG
SSSSR[RR=R:R8NHGRR+L
G;SSSS	RRRRR:=[RR+4S;
SHSSVGRLRI>RH-8L4sRFR8NHGRR>INH8-04RE
CMRRRRRRRRRRRRRHRRVRR[<bRIs08RERCMRRSS-x-RCRsFCCG0MS8
SSSSSl1k)5FI[:2R= RZ)(m4;S
SSCSSMH8RVS;
SSSSH	VRRI<RbRs80MECRSRSRR--xFCsR0CGC
M8SSSSSkS1lI)F5R	2:Z=R 4)m(S;
SSSSCRM8H
V;SSSSCHD#VHRN8<GRR0jRE
CMSSSSSRHV[RR<jER0CRMRSRSS-N-R8#[k0ER0CMRH8COH#FRl8FkDRNIlGS
SSSSS[=R:R+[RRI.*l;NG
SSSSMSC8VRH;S
SSHSSVRR	<RRj0MEC
SSSS	SSRR:=	RR+.l*IN
G;SSSSS8CMR;HV
SSSSVSHR<[RRRLG0MEC
SSSS1SSkFl)I25[RR:=Zm )4
(;RRRRRRRRRRRRRCRRDV#HR<[RRsIb8ER0CRMRR-RR-CRxsCFRGM0C8S
SSSSS1)klF[I52=R:R)Z m;4(
SSSSMSC8VRH;S
SSHSSVRR	<L=RGER0CSM
SSSSSl1k)5FI	:2R= RZ)(m4;R
RRRRRRRRRRRRRR#CDH	VRRI<RbRs80MECRRRRRR--xFCsR0CGC
M8SSSSSkS1lI)F5R	2:Z=R 4)m(S;
SSSSCRM8H
V;SSSSCCD#
SSSSkS1lI)F5R[2:u=RsqF8s$sN58NHGH*I8LL+GR25RvWz-84RF0IMFRRRj
2;RRRRRRRRRRRRRHRRVRR	<bRIs08RE
CMSSSSSkS1lI)F5R	2:u=RsqF8s$sN58NHGH*I8LL+G.25*vWz-84RF0IMFzRWv
2;SSSSS8CMR;HV
SSSS8CMR;HV
SSSCRM8DbFF;-RR-GRL
SSS-O-RFCMPs00RENCRs$sNRRFVOMEk	H#RMR0FNNMRs$sNRRFVL#H0
RRRRRRRRFRVsNRHGMRHR0jRFbRIs48-RFDFbS
SSFSVsGRDRRHMjFR0RvWz-D4RF
FbSSSSSl1k)eFICHO5NWG*zDv+G:2R=kR1lI)F5GHN2G5D2S;
SCSSMD8RF;FbR-R-R
DGSCSSMD8RF;FbR-R-RGHN
SSS-q-R808REsCRF[IRkR#0ONsC0RC800FREsCRkHMMM#oRkRl
RRRRRRRR)1kMk:lR=kR)Ml1kR1+RkFl)IOeC;S
SCRM8DbFF;-RR-xRHGS
S-a-REFCRkk0b0sRbFO8k0#RHRs8CP8HCRFVslER0CkRsMMMHokR#lR
RRRRRu7)mRR<=)1kMkNl5I0H8EI+LHE80-84RF0IMF2Rj;C
SMb8RsCFO#N#R8s8bF
8;
8CMRFLDO;	#
-
-R****************************************************************-RR--
-R-
-R0 MHR0$7DCON0sNHRFMVRFskHM#o8MCRDlk0DHbH
Cs-
-R-a-RERH#H0#RElCRNRHMCHM00V$RF0sREkCRMo#HMRC8l0kDHHbDCRs3RCaERF0IRONsECH0Os0kC-#
-CR8VCHM8CRLDRFIkR#C0RECCHM00#HCRFNLPRC,NRM8l0k#RRLCD0N#RRHM0#EHRDVHCR3Ra
EC-0-RINFRsHOE00COk#sCRCNsRC0ERoDFHPORCHs#FNMRM08RELCRD	FORsPC#MHF3-
-R-
-R****************************************************************-RR-D

HNLssH$RC;CC
Ck#RCHCC03#8F_Do_HO4c4n3DND;#
kCCRHC#C30D8_FOoH_HNs0NE3D
D;kR#CHCCC38#0_oDFHkO_Mo#HM3C8N;DD
H
DLssN$$R#MHbDV
$;kR#C#b$MD$HV30N0skHL03C#N;DD
H
DLssN$sRFO;Nd
Ck#ROFsNFd3sOONF3lbN;DD
M
C0$H0Rpvza#RH
RRRRMoCCOsH5R
RRRRRR8IH0RER:MRH0CCos=R:R;.c
RRRRRRRN8IH0:ERR0HMCsoCRR:=4
.;RRRRRLRRI0H8ERR:HCM0oRCs:4=R.S
SR
2;RRRRb0Fs5S
SRRqRRRR:H#MR0D8_FOoH_OPC05FsN8IH0-ER4FR8IFM0R;j2
RSSARRRRH:RM0R#8F_Do_HOP0COFLs5I0H8E4R-RI8FMR0Fj
2;SuSR)Rm7:kRF00R#8F_Do_HOP0COFIs5HE80RR-48MFI0jFR2R
RRRRRR
2;RNRR0H0sLCk0Rs\3N\M	RH:RMo0CC
s;RNRR0H0sLCk0Rl\3FD8kC:\RRs#0H;Mo
RRRNs00H0LkC3R\bCF8l:\RR0HMCsoC;R
RR0N0skHL0\CR38bFCklL#:\RRs#0H;Mo
RRRNs00H0LkC3R\C_M80CsC\RR:HCM0o;Cs
RRRNs00H0LkC3R\LHCoMs_0CRC\:MRH0CCosR;
R0RN0LsHkR0C\C3slCFP__MFIMNs\RR:HCM0o;Cs
8CMRpvza
;
-*-R*************************************************************R**R
---
-R-D-RFOoHRONsECH0Os0kCV#RFmsRsRON6-
-R-
-R****************************************************************-RR-N

sHOE00COkRsCDHFoOVRFRpvza#RH
-
-RMVH8ER0CNRDssoCR8IH05ERI0H8EFNRsHRI8L0E2R

RkRVMHO0F#MRkIb5HE80NI,RHE80LRR:HCM0o2CsR0sCkRsMHCM0oRCsHR#
RCRLo
HMRRRRRVRHRH5I8N0ERI>RHE80L02RE
CMRRRRRRRRR0sCkRsMI0H8E
N;RRRRRDRC#RC
RRRRRRRRskC0sIMRHE80LR;
RRRRR8CMR;HV
RRRCRM8#;kb
-
-RMVH8ER0ClR#NCDDsHRI8R0E58IH0RENFIsRHE80L
2
RVRRk0MOHRFMH5MVI0H8ERN,I0H8E:LRR0HMCsoC2CRs0MksR0HMCsoCR
H#RLRRCMoH
RRRRHRRVIR5HE80NRR<I0H8ERL20MEC
RRRRRRRRCRs0MksR8IH0;EN
RRRRCRRD
#CRRRRRRRRR0sCkRsMI0H8E
L;RRRRRMRC8VRH;R
RR8CMRVHM;-

-ER0CFRVDIDFHRMoCkM#sRC#00ENR8IH0REAHN#RD$IN#sRoCCN0sER0NFMRsJRCkRND0IFRHE80q-
-RHk#M'oR#'kbR8NMRM'HV
'3
RRRO#FM00NMR8IH0REq:MRH0CCos=R:RVHM5HNI8,0ERHLI820E;R
RRMOF#M0N0HRI8A0ERH:RMo0CC:sR=kR#bI5NHE80,IRLHE802
;
-0-REOCRFFlbM0CMRswH#s0uFO8k05#R#RCCNPLFC
2
RORRFFlbM0CMRswH#s0uFO8k0R#
RCRoMHCsOR5
RRRRR8IH0REq:MRH0CCosR;
RRRRR8IH0REA:MRH0CCosR
RR
2;RbRRFRs05R
RRRRRq:RRRRHMR8#0_oDFHPO_CFO0sI5NHE80-84RF0IMF2Rj;R
RRRRRA:RRRRHMR8#0_oDFHPO_CFO0sI5LHE80-84RF0IMF2Rj;R
RRRRRq:ARR0FkR8#0_oDFHPO_CFO0sI5LHE80*HNI8-0E4FR8IFM0R
j2RRRRR-R-R*ARRRq
R;R2
RRRCRM8ObFlFMMC0
;
-0-REOCRFFlbM0CMR8N8CssaC5CR#RCCNPLFC
2
RORRFFlbM0CMR8N8CssaCRC
RCRoMHCsOR5
RRRRR8IH0REq:MRH0CCosR;
RRRRR8IH0REA:MRH0CCosR
RR
2;RbRRFRs05R
RRRRRqRARRRRR:MRHR8#0_oDFHPO_CFO0sI5LHE80*HNI8-0E4FR8IFM0R;j2
RRRRbRRskF8O:0RR0FkR8#0_oDFHPO_CFO0sI5LHE80+HNI8-0E4FR8IFM0R
j2RRRRR-R-R*ARRRq
R;R2
RRRCRM8ObFlFMMC0
;
R#RRHNoMD_RNNRkGR#:R0D8_FOoH_OPC05FsI0H8E4q-RI8FMR0Fj
2;R#RRHNoMD_RLNRkGR#:R0D8_FOoH_OPC05FsI0H8E4A-RI8FMR0Fj
2;R#RRHNoMDLRNRRRRR#:R0D8_FOoH_OPC05FsN8IH0LE*I0H8ER-48MFI0jFR2R;
RHR#oDMNR#sCkRD0:0R#8F_Do_HOP0COFNs5I0H8EI+LHE80-84RF0IMF2Rj;-

-ER0CHRVsR#0NEsOHO0C0CksRsVFRC0ERDlk0DHb$RR-NNMRs$sNR#LNCl8RkHD0bCDHsL

CMoHRR
RRR--1bINRNqRMA8RRRHVMCCO#s#N$
3RRHRRVNqDssoCAH:RVNR5I0H8ERR>L8IH0RE2oCCMsCN0
RRRRVRRFFsDF:b.RsVFRHHRMRRj0LFRI0H8ER-4oCCMsCN0
RRRRRRRR0RN0LsHkR0C\N3sMR	\FsVRCqo#RD:RNDLCRRH#jS;
S0SN0LsHkR0C\C3slCFP__MFIMNs\VRFRosC#:qRRLDNCHDR#;R4
RRRRRRRR0RN0LsHkR0C\N3sMR	\FsVRCAo#RD:RNDLCRRH#jS;
S0SN0LsHkR0C\C3slCFP__MFIMNs\VRFRosC#:ARRLDNCHDR#;R4
RRRRLRRCMoH
RRRRRRRRCRso:#qRHRbbkCLVR
RRRRRRbRRFRs0l5Nb
RRRRRRRRRRRR=QR>5RAH
2,RRRRRRRRRRRRm>R=RNN_kHG52R
RRRRRR2RR;R
RRRRRRsRRCAo#:bRRHLbCkRV
RRRRRRRRb0FsRblN5R
RRRRRRRRRRRRQ=q>R5,H2
RRRRRRRRRRRR=mR>_RLN5kGHR2
RRRRRRRR2R;
RRRRR8CMRMoCC0sNCFRVsFDFb
.;
RRRRVRRFFsDF:b4RsVFRHHRMIRLHE80RR0FN8IH04E-RMoCC0sNCR
RRRRRRNRR0H0sLCk0Rs\3N\M	RRFVs#CoARR:DCNLD#RHR
j;SNSS0H0sLCk0Rs\3CPlFCF_M_sINMF\RVCRsoR#A:NRDLRCDH4#R;R
RRRRRLHCoMR
RRRRRRsRRCAo#:bRRHLbCkRV
RRRRRRRRb0FsRblN5R
RRRRRRRRRRRRQ=q>R5,H2
RRRRRRRRRRRR=mR>_RLN5kGHR2
RRRRRRRR2R;
RRRRR8CMRMoCC0sNCFRVsFDFb
4;RCRRMo8RCsMCNR0CHDVqNCsos
A;
RRR-z-R#qCRRA&RR0IHE0FkRN#IbMbHoR3
RVRHqN#lDsDCAH:RVNR5I0H8E=R<RHLI820ERMoCC0sNCR
RRRRRVDFsFNFb:FRVsRRHHjMRRR0FN8IH04E-RMoCC0sNCR
RRRRRRNRR0H0sLCk0Rs\3N\M	RRFVs#CoBRR:DCNLD#RHR
j;SNSS0H0sLCk0Rs\3CPlFCF_M_sINMF\RVCRsoR#B:NRDLRCDH4#R;R
RRRRRRNRR0H0sLCk0Rs\3N\M	RRFVs#Co1RR:DCNLD#RHR
j;SNSS0H0sLCk0Rs\3CPlFCF_M_sINMF\RVCRsoR#1:NRDLRCDH4#R;R
RRRRRLHCoMR
RRRRRRsRRCBo#:bRRHLbCkRV
RRRRRRRRb0FsRblN5R
RRRRRRRRRRRRQ=q>R5,H2
RRRRRRRRRRRR=mR>_RNN5kGHR2
RRRRRRRR2R;
RRRRRRRRs#Co1R:RbCHbL
kVRRRRRRRRRsbF0NRlbR5
RRRRRRRRRQRRRR=>A25H,R
RRRRRRRRRRRRm=L>R_GNk5
H2RRRRRRRRR
2;RRRRRMRC8CRoMNCs0VCRFFsDF;bN
R
RRRRRVDFsFLFb:FRVsRRHHNMRI0H8EFR0RHLI8-0E4CRoMNCs0RC
RRRRRRRRNs00H0LkC3R\s	NM\VRFRosC#:7RRLDNCHDR#;Rj
SSSNs00H0LkC3R\sFClPMC_FN_IsRM\FsVRC7o#RD:RNDLCRRH#4R;
RRRRRoLCHRM
RRRRRRRRs#Co7R:RbCHbL
kVRRRRRRRRRsbF0NRlbR5
RRRRRRRRRQRRRR=>A25H,R
RRRRRRRRRRRRm=L>R_GNk5
H2RRRRRRRRR
2;RRRRRMRC8CRoMNCs0VCRFFsDF;bL
RRRCRM8oCCMsCN0RqHV#DlNDACs;R

RHRws1#00:CbRswH#s0uFO8k0R#
RRRRRMoCCOsHRblNRR5
RRRRRRRRI0H8E=qR>HRI8q0E,R
RRRRRRIRRHE80A>R=R8IH0
EARRRRR
R2RRRRRFRbsl0RN5bR
RRRRRRRRRRq=N>R_GNk,R
RRRRRRARRRR=>Lk_NGR,
RRRRRRRRq=AR>LRN
RRRR2RR;R

R8Rq8aCss.CCRN:R8s8CaCsC
RRRRoRRCsMCHlORN5bR
RRRRRRRRHRI8q0ERR=>I0H8E
q,RRRRRRRRR8IH0REA=I>RHE80AR
RRRRR2R
RRRRRb0FsRblNRR5
RRRRRRRRq=AR>LRN,R
RRRRRRbRRskF8O=0R>CRs#0kD
RRRR2RR;R

RuRR)Rm7<s=RCD#k0H5I8-0E4FR8IFM0R;j2
8CMRoDFH
O;
R--****************************************************************R-R-
R--
R--LODF	k_lDN0RsHOE00COk#sCRsVFROmsN
R6-
-R-*-R*************************************************************R**R
--
ONsECH0Os0kCDRLF_O	l0kDRRFVvazpR
H#
-S-RsbkbCF#:CRs0Mks#ER0CCRMIHRI8R0ELCN#8MRFROCGCR##L#H0RHLCMboRsCC#MR0
RkRVMHO0FbMRNW##HE80RR5
RRRRRMOF#M0N0FRl88IH0:ERR0HMCsoC;R
RRRRRO#FM00NMR8FDW0H8ERR:HCM0o2Cs
sSSCs0kMMRH0CCos#RH
CSLoRHMRR--b#N#W0H8ER
RRRRRHlVRFH8I8R0E>RR.0MECR-R-R#lF0NR0	0CRERH#LMsNOSE
SCSs0MksR8FDW0H8ES;
S#CDHlVRFH8I8R0E=RR.0MEC
SSSskC0sFMRDH8W8-0E.S;
S#CDHlVRFH8I8R0E=RR40MEC
SSSskC0sFMRDH8W8-0E4S;
S#CDHlVRFH8I8R0E=RRj0MEC
SSSskC0sFMRDH8W8;0E
CSSDR#CRSSSS-SR-ER0HH#R#kR#bVCsDkkF#S
SS0sCkRsMFWD8HE80;S
SCRM8H
V;S8CMR#bN#8WH0
E;
-S-RsbkbCF#:CRs0Mks#RR4HMVRCRC808FRFHRbbHCDMoHM
kSVMHO0FNMRM$ND#HC_M0bk_8IH0NE5I,H8RHLI8RR:HCM0o2CsR0sCkRsMHCM0oRCsHS#
LHCoMS
SH5VR5HNI8RR>4R(2NRM85HLI8RR>42(2RC0EMS
SS0sCkRsM4R;
RRRRR8CMR;HV
sSSCs0kM;Rj
MSC8MRNN#D$CM_Hb_k0I0H8E
;
R-RR-HRVM08RE#CRlDNDCIsRHE80RH5I8R0EFNsRI0H8ER2
RkRVMHO0FHMRMIV5HE80,IRNHE80RH:RMo0CCRs2skC0sHMRMo0CCHsR#R
RRoLCHRM
RRRRRRHV58IH0<ERRHNI820ERC0EMR
RRRRRRsRRCs0kMHRI8;0E
RRRRCRRD
#CRRRRRRRRR0sCkRsMN8IH0
E;RRRRRMRC8VRH;R
RR8CMRVHM;R

RFROMN#0MW0RzRvRRRR:HCM0oRCs:4=R(S;
SSSSSRR
RFROMN#0MN0RICH8RRR:HCM0oRCs:H=RMIV5HE80,IRNHE802S;
O#FM00NMRHLI8RCR:MRH0CCos=R:RVHM58IH0RE,L8IH0;E2
SSSSRSS
RRRO#FM00NMRFNl8RRR:MRH0CCos=R:RHNI85C-5N55ICH8+vWz-/42W2zv-*42W2zv;R
RRMOF#M0N0lRLFR8RRH:RMo0CC:sR=IRLH-8C5555L8IHCz+Wv2-4/vWz22-4*vWz2S;
SSSSSRR
RFROMN#0MN0RIRH8SRR:HCM0oRCs:b=RNW##HE805FNl8N,RICH82R;
RFROMN#0ML0RIRH8SRR:HCM0oRCs:b=RNW##HE805FLl8L,RICH82
;
RORRF0M#NRM0M8CC_bbHCMDHCRR:HCM0oRCs:N=RM$ND#HC_M0bk_8IH0NE5I0H8EL,RI0H8E
2;SSSSSSRRR#
SHNoMD4RCRRRRR:SRR8#0_oDFHPO_CFO0sR548MFI0jFR2S;
#MHoNCDR.RRRRRRS:0R#8F_Do_HOP0COF4s5RI8FMR0Fj
2;SSSSSSRRRR
RRo#HMRNDqH0slRRRR#:R0D8_FOoH_OPC05FsN8IHCR-48MFI0jFR2R;
RHR#oDMNRsA0HRlRRRR:#_08DHFoOC_POs0F5HLI84C-RI8FMR0Fj
2;
RRR#MHoNqDRblsHCRRR:0R#8F_Do_HOP0COFNs5I-H84FR8IFM0R;j2
RRR#MHoNADRblsHCRRR:0R#8F_Do_HOP0COFLs5I-H84FR8IFM0R;j2
RRR#MHoN1DRE0FsuRRR:0R#8F_Do_HOP0COFNs5I+H8L8IH-84RF0IMF2Rj;S
SSSSSRR
RRo#HMRND)kC#DR04R#:R0D8_FOoH_OPC05FsN8IHCI+LH-8C4FR8IFM0R;j2
RRR#MHoN)DRCD#k0RGR:0R#8F_Do_HOP0COFNs5ICH8+HLI84C-RI8FMR0Fj
2;R#RRHNoMDCR)#0kDN:RRR8#0_oDFHPO_CFO0sI5NH+8CL8IHCR-48MFI0jFR2R;
RHR#oDMNR#)CkLD0RRR:#_08DHFoOC_POs0F5HNI8LC+ICH8-84RF0IMF2Rj;R
RRo#HMRND)kC#DR0CR#:R0D8_FOoH_OPC05FsN8IHCI+LH-8C4FR8IFM0RRj2:5=RFC0Es=#R>jR''
2;
RRR#MHoNuDRs4F8_GNk,sRuF_84sRC#RRR:#_08DHFoOC_POs0F5HNI8LC+ICH8-84RF0IMF2Rj;R
RRo#HMRNDu8sF4RRRR#:R0D8_FOoH_OPC05FsN8IHCI+LH-8C4FR8IFM0R;j2
RRR#MHoNuDRs.F8RRRR:0R#8F_Do_HOP0COFIs5HE80-84RF0IMF2Rj;S

ObFlFMMC0.ReABpmiS
SoCCMsRHO5S
SSHNI8R0E:MRH0CCos=R:RHNI8S;
SISLHE80RH:RMo0CC:sR=IRLH
8;SMSSC_C8bCHbDCHMRH:RMo0CC:sR=CRMCb8_HDbCH2MC;S
Sb0FsRS5
SRSqR:RRRRHMR8#0_oDFHPO_CFO0sI5NH48-RI8FMR0Fj
2;SASSRRRR:MRHR0R#8F_Do_HOP0COFLs5I-H84FR8IFM0R;j2
SSSu7)mRF:Rk#0R0D8_FOoH_OPC05FsN8IH+HLI8R-48MFI0jFR2
2;S8CMRlOFbCFMM
0;
oLCHRMR-L-RD	FO_Dlk0S

-b-RkFsb#RC:0CN	RsONCVRFRC0ERN4RM.8R-0LHR#ONCS#
-0-R$RbCRRR:OLFlH0MNHNFMD-
S-MRHb#k0Rq:R,
RASR--Fbk0k:0#Rmu)7-
S-sR0H0lREHCRM0bk#FR0RRLCMIFRHs8CRN0EMER0CkRF00bk
VSH_MoC:VRHRC5MCb8_HDbCHRMC=2R4RMoCC0sNCS
S0lsHH:0qRsVFRHHRMRRj0NFRICH8-o4RCsMCN
0CSNSS0H0sLCk0Rs\3N\M	RRFVs#CoqRR:DCNLD#RHR
j;SNSS0H0sLCk0Rb\3Fl8C\VRFRosC#:qRRLDNCHDR#;RH
SSSNs00H0LkC3R\bCF8l#Lk\VRFRosC#:qRRLDNCHDR#qR""S;
S0SN0LsHkR0C\F3l8CkD\VRFRosC#:qRRLDNCHDR#vR"z"pa;S
SS0N0skHL0\CR3lsCF_PCMIF_N\sMRRFVs#CoqRR:DCNLD#RHR
4;SCSLo
HMSsSSCqo#:bRRHLbCkSV
SbSSFRs0l5Nb
SSSSRSQ=q>R5,H2
SSSSRSm=q>R0lsH5
H2SSSS2S;
S8CMRMoCC0sNCsR0H0lHq
;
RSRS0lsHH:0ARsVFRHHRMRRj0LFRICH8-o4RCsMCN
0CSNSS0H0sLCk0Rs\3N\M	RRFVs#CoARR:DCNLD#RHR
j;SNSS0H0sLCk0Rb\3Fl8C\VRFRosC#:ARRLDNCHDR#;RH
SSSNs00H0LkC3R\bCF8l#Lk\VRFRosC#:ARRLDNCHDR#AR""S;
S0SN0LsHkR0C\F3l8CkD\VRFRosC#:ARRLDNCHDR#vR"z"pa;S
SS0N0skHL0\CR3lsCF_PCMIF_N\sMRRFVs#CoARR:DCNLD#RHR
4;SCSLo
HMSsSSCAo#:bRRHLbCkSV
SbSSFRs0l5Nb
SSSSRSQ=A>R5,H2
SSSSRSm=A>R0lsH5
H2SSSS2S;
S8CMRMoCC0sNCsR0H0lHAS;
CRM8oCCMsCN0R_HVo;CM
H
SVC_oMRj:H5VRM8CC_bbHCMDHCRR=jo2RCsMCN
0CS0SqsRHl<q=R5HNI84C-RI8FMR0Fj
2;S0SAsRHl<A=R5HLI84C-RI8FMR0Fj
2;S8CMRMoCC0sNCVRH_MoCj
;
SR--sFClP0CRECCRGN0sR0LH#0RNRC0ERAp1R8CM
RRRbMskC:H0RFbsO#C#R05qs,HlRsA0H
l2SoLCHRMR-b-RsCFO#b#RsCkMHS0
SRHVN8lFR4=RRC0EMS
SSRC4<'=Rj&'RRsq0Hjl52S;
SbSqsCHlRR<=qH0slI5NH-8C4FR8IFM0R;42
CSSDV#HRFNl8RR=.ER0CRM
RRRRRRRRC<4R=0Rqs5Hl4FR8IFM0R;j2
SSSqHbsl<CR=0Rqs5HlN8IHCR-48MFI0.FR2R;
RRRRR#CDCS
SSRC4<'=Rj&'RR''j;S
SSsqbHRlC<q=R0lsH;S
SCRM8H
V;
HSSVlRLF=8RR04RE
CMSCSS.=R<R''jRA&R0lsH5;j2
SSSAHbsl<CR=0RAs5HlL8IHCR-48MFI04FR2S;
S#CDHLVRlRF8=RR.0MEC
RRRRRRRR.RCRR<=AH0slR548MFI0jFR2S;
SbSAsCHlRR<=AH0slI5LH-8C4FR8IFM0R;.2
RRRRCRRD
#CSCSS.=R<R''jR'&Rj
';SASSblsHC=R<RsA0H
l;SMSC8VRH;C
SMb8RsCFO#b#RsCkMH
0;
-S-RDvk0DHb$$RLRC0ER0CGsLNRHR0#HIVRCNREPFCRMFCRsIR0FGRC0RsNL#H0RRFVqH
SV4_N:VRHRl5NF=8RRR42oCCMsCN0
HSSV4_NLRj:H5VRL8lFRR<=jsRFRFLl8RR>.o2RCsMCN
0CS)SSCD#k0<NR=mRBh1e_ap7_mBtQ_Be a5m)jN,RICH8+HLI8RC2IMECR45C5Rj2=jR''
2RSSSSSRSRCCD#Ra X5sAbH,lCRHNI8LC+ICH82R;
RRRRR8CMRMoCC0sNCVRH_LN4jS;
S_HVN44L:VRHRl5LF=8RRR42oCCMsCN0
SSS)kC#DR0N<B=Rm_he1_a7pQmtB _eB)am5Rj,N8IHCI+LH28CRCIEMCR5425jR'=RjR'2
SSSSRSSR#CDCXR ab5AsCHlR'&RjR',N8IHCI+LH28C;R
RRRRRCRM8oCCMsCN0R_HVN44L;S
SHNV_4:L.RRHV5FLl8RR=.o2RCsMCN
0CS)SSCD#k0<NR=mRBh1e_ap7_mBtQ_Be a5m)jN,RICH8+HLI8RC2IMECR45C5Rj2=jR''
2RSSSSSRSRCCD#Ra X5sAbHRlC&jR''RR&',j'RHNI8LC+ICH82R;
RRRRR8CMRMoCC0sNCVRH_LN4.S;
CRM8oCCMsCN0R_HVN
4;S_HVNR.:H5VRN8lFR.=R2CRoMNCs0RC
RRRRRo#HMRNDMEF1H,V0RH#EV80C,8RN8RC8:0R#8F_Do_HOP0COFNs5ICH8+HLI84C-RI8FMR0Fj
2;SoLCHSM
S_HVNj.L:VRHRl5LF<8R=RRjFLsRlRF8>2R.RMoCC0sNCR
RRMSSFH1EV<0R=XR ab5AsCHl,IRNH+8CL8IHC
2;RRRRRMRC8CRoMNCs0HCRV._NL
j;SVSH_LN.4H:RVLR5lRF8=2R4RMoCC0sNCR
RRMSSFH1EV<0R=XR ab5AsCHlR'&RjR',N8IHCI+LH28C;R
RRRRRCRM8oCCMsCN0R_HVN4.L;S
SHNV_.:L.RRHV5FLl8RR=.o2RCsMCN
0CRSRRS1MFE0HVRR<= 5XaAHbsl&CRR''jR'&RjR',N8IHCI+LH28C;R
RRRRRCRM8oCCMsCN0R_HVN..L;R
RSES#HCV08=R<R#MFE0HV5HNI8LC+ICH8-8.RF0IMF2RjR'&Rj
';S8SN8RC8R=R<R1MFE0HVR#+RE0HVC
8;RSRR)kC#DR0N<B=Rm_he1_a7pQmtB _eB)am5Nj,ICH8+HLI8RC2IMECR45CR"=Rj2j"
SSSSRSRCCD#R1MFE0HVRCIEMCR54RR=""j42S
SSRSSR#CDCER#HCV08ERIC5MRC=4RRj"4"S2
SSSSRDRC#NCR888C;C
SMo8RCsMCNR0CHNV_.
;
SR--v0kDH$bDRRL$0RECCsG0NHRL0H#RVCRIRPENCMRFCsRFRF0IR0CGsLNRHR0#FAVR
VSH_:L4RRHV5FLl8RR=4o2RCsMCN
0CSVSH_NL4jH:RVNR5lRF8<j=RRRFsN8lFR.>R2CRoMNCs0SC
SCS)#0kDL=R<RhBmea_17m_pt_QBea Bmj)5,IRNH+8CL8IHCI2RERCM55C.j=2RR''j2SR
SSSSSCRRDR#C 5XaqHbslRC,N8IHCI+LH28C;R
RRRRRCRM8oCCMsCN0R_HVLj4N;S
SHLV_4:N4RRHV5FNl8RR=4o2RCsMCN
0CS)SSCD#k0<LR=mRBh1e_ap7_mBtQ_Be a5m)jN,RICH8+HLI8RC2IMECR.5C5Rj2=jR''
2RSSSSSRSRCCD#Ra X5sqbHRlC&jR''N,RICH8+HLI8;C2
RRRRCRRMo8RCsMCNR0CHLV_4;N4
HSSV4_LNR.:H5VRN8lFR.=R2CRoMNCs0SC
SCS)#0kDL=R<RhBmea_17m_pt_QBea Bmj)5,IRNH+8CL8IHCI2RERCM55C.j=2RR''j2SR
SSSSSCRRDR#C 5XaqHbsl&CRR''jR'&RjR',N8IHCI+LH28C;R
RRRRRCRM8oCCMsCN0R_HVL.4N;C
SMo8RCsMCNR0CHLV_4S;
HLV_.H:RVLR5lRF8=2R.RMoCC0sNCR
RRRRR#MHoNMDRFH1EVR0,#VEH0,C8R8N8C:8RR8#0_oDFHPO_CFO0sI5NH+8CL8IHCR-48MFI0jFR2S;
LHCoMS
SHLV_.:NjRRHV5FNl8=R<RFjRslRNF>8RRR.2oCCMsCN0
RRRSFSM1VEH0=R<Ra X5sqbH,lCRHNI8LC+ICH82R;
RRRRR8CMRMoCC0sNCVRH_NL.jS;
S_HVL4.N:VRHRl5NF=8RRR42oCCMsCN0
RRRSFSM1VEH0=R<Ra X5sqbHRlC&jR''N,RICH8+HLI8;C2
RRRRCRRMo8RCsMCNR0CHLV_.;N4
HSSV._LNR.:H5VRN8lFR.=R2CRoMNCs0RC
RSRSMEF1HRV0< =RXqa5blsHCRR&'Rj'&jR''N,RICH8+HLI8;C2
RRRRCRRMo8RCsMCNR0CHLV_.;N.
#SSE0HVC<8R=FRM1VEH0I5NH+8CL8IHCR-.8MFI0jFR2RR&';j'
RRRRNRR888CR<RR=FRM1VEH0RR+#VEH0;C8
)SSCD#k0<LR=mRBh1e_ap7_mBtQ_Be a5m)jN,RICH8+HLI8RC2IMECR.5CR"=Rj2j"
SSSSRSRCCD#R1MFE0HVRCIEMCR5.RR=""j42S
SSRSSR#CDCER#HCV08ERIC5MRC=.RRj"4"S2
SSSSRDRC#NCR888C;C
SMo8RCsMCNR0CHLV_.
;
SR--v0kDH$bDRC0ER0CGsLNRHR0#0CFo0sECRRHVIECRNRPCCsG0NH#RMRRqNRM8AH
SV#_C:VRHRN55l=F84sRFRFNl82=.R8NMRl5LF48=RRFsL8lF=2.2RMoCC0sNCS
S)kC#D50Cd<2R=4RC5R42NRM8Cj452MRN8.RC5R42NRM8Cj.52S;
S#)CkCD05R.2<5=RC4452MRN8MR5FC0R425j2MRN8.RC5242R
FsSSSSSRSR55C44N2RMC8R.254R8NMRF5M0.RC52j22S;
S#)CkCD05R42<5=RC4452MRN8MR5FC0R.2542MRN8.RC52j2R
FsSSSSSRSR55C44N2RM58RMRF0Cj452N2RMC8R.25j2sRF
SSSSRSSRM55FC0R42542MRN84RC5Rj2NRM8C4.52F2RsS
SSSSSRCR5425jR8NMR5C.4N2RM58RMRF0Cj.52;22
)SSCD#k0jC52=R<R5C4jN2RMC8R.25j;S
SHsV_C:#CRRHV5HNI8LC+ICH8Rc>R2CRoMNCs0SC
SCS)#0kDCI5NHR8C+IRLHR8C-RR48MFI0cFR2=R<RhBmea_17m_pt_QBea Bmj)5,IRNH+8CL8IHCcR-2S;
S8CMRMoCC0sNCVRH_#sCCS;
CRM8oCCMsCN0R_HVC
#;
lSLk:D0RRHVN8IHCRR>.MRN8IRLHR8C>RR.oCCMsCN0
lSSkGD0GRR:ep.Am
BiSoSSCsMCHlORN5bR
SSSSNSSI0H8E>R=RHNI8S,
SSSSSHLI8R0E=L>RI,H8
SSSSMSSC_C8bCHbDCHMRR=>M8CC_bbHCMDHCS2
SFSbsl0RN5bR
SSSSRSqR=RR>bRqsCHl,S
SSASSRRRR=A>RblsHCS,
SSSSu7)mRR=>1sEF0;u2
MSC8CRoMNCs0LCRl0kD;S

CCG0M08H:sRbF#OC#1R5E0FsuS2
LHCoM-RR-sRbF#OC#GRC08CMHS0
S#)Ck4D0RR<= 5Xa1sEF0Ru,N8IHCI+LH28C;C
SMb8RsCFO#C#RGM0C8;H0
N
SL8lFjH:RVNR5l>F8.sRFRFNl82=jR8NMRl5LF.8>RRFsL8lF=Rj2oCCMsCN0
)SSCD#k0<GR=CR)#0kD4S;
CRM8oCCMsCN0RlNLF;8j
R
RSlNLF:84RRHV5FNl8R=4NRM85FLl8R>.FLsRl=F8jR22F5sR5FNl8R>.FNsRl=F8jN2RML8Rl=F84o2RCsMCN
0CSCS)#0kDG=R<R#)Ck4D05HNI8LC+ICH8-8.RF0IMF2RjR'&Rj
';S8CMRMoCC0sNCLRNl4F8;S

NFLl8R.:H5VRN8lF=N4RML8Rl=F84F2RsNR5l=F8.MRN8LR5l>F8.sRFRFLl82=j2sRFRN55l>F8.sRFRFNl82=jR8NMRFLl82=.RMoCC0sNCS
S)kC#DR0G<)=RCD#k0N45ICH8+HLI8dC-RI8FMR0Fj&2RRj"j"S;
CRM8oCCMsCN0RlNLF;8.
N
SL8lFdH:RVNR5l=F8.MRN8lRLF48=2sRFRl5NF48=R8NMRFLl82=.RMoCC0sNCS
S)kC#DR0G<)=RCD#k0N45ICH8+HLI8cC-RI8FMR0Fj&2RRj"jj
";S8CMRMoCC0sNCLRNldF8;R

RLSNlcF8:VRHRl5NF.8=R8NMRFLl82=.RMoCC0sNCS
S)kC#DR0G<)=RCD#k0N45ICH8+HLI86C-RI8FMR0Fj&2RRj"jj;j"
MSC8CRoMNCs0NCRL8lFc
;
S_HVoCCMsCN0:VRHR555N8lFRj>R2MRN8NR5lRF8<2Rd2sRFRL55lRF8>2RjR8NMRl5LF<8RR2d22CRoMNCs0SC
LHCoMS
SH#V_0CN04H:RV5R5N8lFRj>R2MRN8NR5lRF8<2RdR8NMRl5LF>8RRRj2NRM85FLl8RR<dR22oCCMsCN0
SSSu8sF4k_NG=R<RCR)#0kDNRR+)kC#DR0L+CR)#0kDCS;
S8CMRMoCC0sNCVRH_N#00;C4
HSSV0_#N.0C:VRHRN55lRF8>2RjR8NMRl5NF<8RRRd2NRM85l5LF>8RRR.2F5sRL8lFRj=R2R22oCCMsCN0
SSSu8sF4k_NG=R<RCR)#0kDNS;
S8CMRMoCC0sNCVRH_N#00;C.
HSSV0_#Nd0C:VRHRL55lRF8>2RjR8NMRl5LF<8RRRd2NRM85l5NF>8RRR.2F5sRN8lFRj=R2R22oCCMsCN0
SSSu8sF4k_NG=R<RCR)#0kDLS;
S8CMRMoCC0sNCVRH_N#00;Cd
S
SHbV_H:b4RRHV5CMC8H_bbHCDM=CRRR42oCCMsCN0
SSSLFkVkk0b0V:RFHsRRRHMjFR0RHNI8R0E+IRLHE80-o4RCsMCN
0CSSSSNs00H0LkC3R\s	NM\VRFRosC#:1RRLDNCHDR#;R4
SSSS0N0skHL0\CR3oLCH0M_s\CCRRFVs#Co1RR:DCNLD#RHR
4;SSSSNs00H0LkC3R\sFClPMC_FN_IsRM\FsVRC1o#RD:RNDLCRRH#4S;
SCSLo
HMSSSSs#Co1R:RbCHbL
kVSSSSb0FsRblN5S
SSSSSQ>R=RFus8N4_kHG52S,
SSSSS=mR>sRuF_84s5C#HS2
SSSSS
2;SCSSMo8RCsMCNR0CLFkVkk0b0S;
S8CMRMoCC0sNCVRH_bbH4S;
S_HVbjHb:VRHRC5MCb8_HDbCHRMC=2RjRMoCC0sNCS
SSFus8s4_CN#5I0H8ERR+L8IH0-ERR84RF0IMF2RjRR<=
SSSSFus8N4_kNG5I0H8ERR+L8IH0-ERR84RF0IMF2Rj;SR
S8CMRMoCC0sNCVRH_bbHj
;
SsSuFR84<)=RCD#k0+GRRFus8s4_C
#;S8CMRMoCC0sNCVRH_MoCC0sNC
;
S_HVoCCMsCN0_R4:H5VR5FNl8RR>.N2RM58RL8lFR.>R2o2RCsMCN
0CSsSuFR84<)=RCD#k0
G;S8CMRMoCC0sNCVRH_MoCC0sNC;_4


RS0CGCbM8s:F8RFbsO#C#Rs5uF284
CSLoRHMRR--bOsFCR##CCG0Ms8bFS8
SRHVI0H8ERR>N8IHCRR+L8IHCER0CSM
SsSuFR8.< =RXua5s4F8,HRI820E;S
SCCD#
SSSu8sF.=R<RFus8I45HE80-84RF0IMF2Rj;S
SCRM8H
V;S8CMRFbsO#C#R0CGCbM8s;F8
H
SVH_bb:N4RRHV5CMC8H_bbHCDM=CRRR42oCCMsCN0
LSSkkVF00bk:FRVsRRHHjMRRR0FI0H8ER-4oCCMsCN0
SSSNs00H0LkC3R\s	NM\VRFRosC#:1RRLDNCHDR#;R.
SSSNs00H0LkC3R\C_M80CsC\VRFRosC#:1RRLDNCHDR#;R.
SSSNs00H0LkC3R\bCF8lF\RVCRsoR#1:NRDLRCDHH#R;S
SS0N0skHL0\CR38bFCklL#F\RVCRsoR#1:NRDLRCDH"#Ru7)m"S;
S0SN0LsHkR0C\C3slCFP__MFIMNs\VRFRosC#:1RRLDNCHDR#;R4
LSSCMoH
SSSs#Co1R:RbCHbL
kVSSSSb0FsRblN5S
SSSSSQ>R=RFus8H.52S,
SSSSS=mR>)RumH752S
SS;S2
CSSMo8RCsMCNR0CLFkVkk0b0S;
CRM8oCCMsCN0R_HVbNHb4S;
HbV_HjbN:VRHRC5MCb8_HDbCHRMC=2RjRMoCC0sNCS
Su7)mRR<=u8sF.H5I8-0E4FR8IFM0R;j2
MSC8CRoMNCs0HCRVH_bb;Nj
M
C8DRLF_O	l0kD;



