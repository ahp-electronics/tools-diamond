-- $Header: //synplicity/map202003lat/mappers/lattice/lib/gen_lava1/add.vhd#1 $
@ER--q
77DsHLNRs$Q   ;#
kC RQ # 30D8_FOoH_n44cD3ND
;
b	NONRoCN0sHEH_DL#RH
0RR$RbC#CbC8ba$C#RHRD5#FRI,lHC8kRl,V0N#2C;
MN8RsEH0_LDH;



LDHs$NsR Q  k;
#QCR 3  #_08DHFoO4_4nNc3D
D;kR#CI	Fs3HNs0DE_HNL3D
D;
0CMHR0$qR77H
#
oCCMs5HOI0H8ERR:HCM0o:Cs=U4.R#;Rb8CCR#:Rb8CCaC$bRR:=V0N#R
2;
sbF0
5
qR,A:MRHR8#0_oDFHPO_CFO0sH5I8-0E4FR8IFM0R;j2
R
RRRRRRQRBhH:RM0R#8F_Do;HO
R
m:kRF00R#8F_Do_HOP0COFIs5HE80-84RF0IMF2Rj;B

mRza:kRF00R#8F_Do
HO

2;
8CMR7q7;N

sHOE00COkRsCV0N#RRFVqR77H
#
ObFlFMMC0BRBz7_q7R
RRsbF0R5
RRRRRRqjRRRRRRRRRRRRRRRRRRRRRRRRRRRR:HRRMRRRR71a_tpmQ
B;RRRRRjRARRRRRRRRRRRRRRRRRRRRRRRRRRRRRR:RHRMRRaR17m_pt;QB
RRRRBRRQRhRRRRRRRRRRRRRRRRRRRRRRRRRRRR:RRHMR1RRap7_mBtQ;R
RRRRR1RjRRRRRRRRRRRRRRRRRRRRRRRRRR:RRRkRF0RRR1_a7pQmtBR;
RRRRRzBmaRRRRRRRRRRRRRRRRRRRRRRRRRRR:FRRkR0RR71a_tpmQ;B2
8CMRlOFbCFMM
0;
o#HMRNDOsNs$RRR:0R#8F_Do_HOP0COFRs5I0H8ER-48MFI0jFRR
2;#MHoNODRF0M#_:4RR8#0_oDFH
O;
oLCHSM
zR4:B_BzqR77uam)Ruvq55RqjR2,A25j,QRBhm,R5,j2RsONsj$52
2;RRRRRRRRpR.:VRFsHMRHR04RFHRI8-0E4CRoMNCs0RC
RRRRRRRRRRRRRzRR.RR:B_BzqR77uam)Ruvq55RqHR2,A25H,NROs5s$H2-4,5RmHR2,OsNs$25H2R;
RRRRRCRRMo8RCsMCN;0C
RRRRRRRRzBma=R<RsONsR$5I0H8ER-42
;

8CMR#VN0
;

ONsECH0Os0kCCRl8lHkRRFVqR77H
#
ObFlFMMC0BRBz7_q7R
RRsbF0R5
RRRRRRqjRRRRRRRRRRRRRRRRRRRRRRRRRRRR:HRRMRRRR71a_tpmQ
B;RRRRRjRARRRRRRRRRRRRRRRRRRRRRRRRRRRRRR:RHRMRRaR17m_pt;QB
RRRRBRRQRhRRRRRRRRRRRRRRRRRRRRRRRRRRRR:RRHMR1RRap7_mBtQ;R
RRRRR1RjRRRRRRRRRRRRRRRRRRRRRRRRRR:RRRkRF0RRR1_a7pQmtBR;
RRRRRzBmaRRRRRRRRRRRRRRRRRRRRRRRRRRR:FRRkR0RR71a_tpmQ;B2
8CMRlOFbCFMM
0;
o#HMRNDOsNs$RRR:0R#8F_Do_HOP0COFRs5I0H8ER-48MFI0jFRR
2;#MHoNODRF0M#_:4RR8#0_oDFH
O;
oLCHSM
zR4:B_BzqR77uam)Ruvq55RqjR2,A25j,QRBhm,R5,j2RsONsj$52
2;RRRRRRRRpR.:VRFsHMRHR04RFHRI8-0E4CRoMNCs0RC
RRRRRRRRRRRRRzRR.RR:B_BzqR77uam)Ruvq55RqHR2,A25H,NROs5s$H2-4,5RmHR2,OsNs$25H2R;
RRRRRCRRMo8RCsMCN;0C
RRRRRRRRzBma=R<RsONsR$5I0H8ER-42
;

8CMR8lCH;kl
ONsECH0Os0kCDR#FFIRV7Rq7#RH
F
OlMbFCRM0B_Bzq
77RbRRF5s0
RRRRqRRjRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR:RRHMR1RRap7_mBtQ;R
RRRRRARjRRRRRRRRRRRRRRRRRRRRRRRRRR:RRRMRHRRRR1_a7pQmtBR;
RRRRRhBQRRRRRRRRRRRRRRRRRRRRRRRRRRRR:HRRMRRRR71a_tpmQ
B;RRRRRjR1RRRRRRRRRRRRRRRRRRRRRRRRRRRRRR:RFRk0RaR17m_pt;QB
RRRRBRRmRzaRRRRRRRRRRRRRRRRRRRRRRRRRRR:R0FkR1RRap7_mBtQ2C;
MO8RFFlbM0CM;#

HNoMDNROsRs$RRR:#_08DHFoOC_POs0F5HRI8-0E4FR8IFM0R2jR;H
#oDMNRMOF#40_R#:R0D8_FOoH;L

CMoH
4Sz:BRBz7_q7mRu)vaRqRu5q25j,5RAjR2,B,QhRjm52O,RN$ss52j2;R
RRRRRR.Rp:FRVsRRHH4MRRR0FI0H8ER-4oCCMsCN0
RRRRRRRRRRRRRRRRRz.:BRBz7_q7mRu)vaRqRu5q25H,5RAHR2,OsNs$-5H4R2,m25H,NROs5s$H;22
RRRRRRRR8CMRMoCC0sNCR;
RRRRRBRRmRza<O=RN$ss5HRI8-0E4;R2
C

M#8RD;FI
