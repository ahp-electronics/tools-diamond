library verilog;
use verilog.vl_types.all;
entity i2cfifo_snow_wrap is
    port(
        ack_o           : out    vl_logic;
        dat_o           : out    vl_logic_vector(9 downto 0);
        i2c_tiehi       : out    vl_logic;
        i2c_tielo       : out    vl_logic;
        i2c_wkup        : out    vl_logic;
        irq             : out    vl_logic;
        mrdcmpl         : out    vl_logic;
        pmu_wkup        : out    vl_logic;
        rxfifo_af       : out    vl_logic;
        rxfifo_e        : out    vl_logic;
        rxfifo_f        : out    vl_logic;
        scl_oe_n        : out    vl_logic;
        scl_out         : out    vl_logic;
        sda_oe_n        : out    vl_logic;
        sda_out         : out    vl_logic;
        srdwr           : out    vl_logic;
        txfifo_ae       : out    vl_logic;
        txfifo_e        : out    vl_logic;
        txfifo_f        : out    vl_logic;
        ADDR_LSB_USR    : in     vl_logic_vector(1 downto 0);
        adr_i           : in     vl_logic_vector(3 downto 0);
        alt_scl_in      : in     vl_logic;
        alt_sda_in      : in     vl_logic;
        cfg_sbi_seln    : in     vl_logic;
        clk_cib         : in     vl_logic;
        cs_i            : in     vl_logic;
        dat_i           : in     vl_logic_vector(9 downto 0);
        fifo_rst        : in     vl_logic;
        mc1_mstr_sleep_rx: in     vl_logic;
        mc1_scl_alt_sel : in     vl_logic;
        mc1_sda_alt_sel : in     vl_logic;
        mc1_sda_i_del   : in     vl_logic;
        mc1_sda_o_del   : in     vl_logic;
        por_n           : in     vl_logic;
        presleep_n      : in     vl_logic;
        presleep_n_ctrl_oe: in     vl_logic;
        presleep_n_ctrl_out: in     vl_logic;
        sbi_init_adr    : in     vl_logic_vector(3 downto 0);
        sbi_init_clk    : in     vl_logic;
        sbi_init_cs     : in     vl_logic;
        sbi_init_dat_i  : in     vl_logic_vector(9 downto 0);
        sbi_init_stb    : in     vl_logic;
        sbi_init_we     : in     vl_logic;
        scl_in          : in     vl_logic;
        sda_in          : in     vl_logic;
        sleep_clk       : in     vl_logic;
        stb_i           : in     vl_logic;
        stop_n          : in     vl_logic;
        vcc             : in     vl_logic;
        vss             : in     vl_logic;
        we_i            : in     vl_logic
    );
end i2cfifo_snow_wrap;
