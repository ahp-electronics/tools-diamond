library verilog;
use verilog.vl_types.all;
entity LSC_OR2 is
    port(
        X               : out    vl_logic;
        A1              : in     vl_logic;
        A2              : in     vl_logic;
        VDD             : in     vl_logic;
        VSS             : in     vl_logic;
        VBP             : in     vl_logic;
        VBN             : in     vl_logic
    );
end LSC_OR2;
