library verilog;
use verilog.vl_types.all;
entity char_test_logic is
    port(
        char_out        : out    vl_logic_vector(21 downto 0);
        test_mode       : out    vl_logic_vector(2 downto 0);
        serdes_char_out : out    vl_logic_vector(21 downto 0);
        tck_fleximac    : out    vl_logic;
        char_td         : out    vl_logic_vector(9 downto 0);
        scan_mode       : out    vl_logic;
        scan_in_tx      : out    vl_logic;
        scan_in_rx      : out    vl_logic;
        scan_enable     : out    vl_logic;
        scan_rstn       : out    vl_logic;
        testclk         : out    vl_logic;
        bist_rstn       : out    vl_logic;
        do_bist         : out    vl_logic;
        cptdr           : out    vl_logic;
        shdr            : out    vl_logic;
        bistrtcntdone   : out    vl_logic;
        char_in         : in     vl_logic_vector(12 downto 0);
        char_mode       : in     vl_logic;
        serdes_char_out_prev: in     vl_logic_vector(21 downto 0);
        tck_fleximac_sel: in     vl_logic;
        tck_fleximac_prev: in     vl_logic;
        rd0             : in     vl_logic_vector(9 downto 0);
        rck0            : in     vl_logic;
        tck0            : in     vl_logic;
        rlol0           : in     vl_logic;
        rlos_hi0        : in     vl_logic;
        rlos_lo0        : in     vl_logic;
        pci_connect0    : in     vl_logic;
        pci_det_done0   : in     vl_logic;
        rd1             : in     vl_logic_vector(9 downto 0);
        rck1            : in     vl_logic;
        tck1            : in     vl_logic;
        rlol1           : in     vl_logic;
        rlos_hi1        : in     vl_logic;
        rlos_lo1        : in     vl_logic;
        pci_connect1    : in     vl_logic;
        pci_det_done1   : in     vl_logic;
        rd2             : in     vl_logic_vector(9 downto 0);
        rck2            : in     vl_logic;
        tck2            : in     vl_logic;
        rlol2           : in     vl_logic;
        rlos_hi2        : in     vl_logic;
        rlos_lo2        : in     vl_logic;
        pci_connect2    : in     vl_logic;
        pci_det_done2   : in     vl_logic;
        rd3             : in     vl_logic_vector(9 downto 0);
        rck3            : in     vl_logic;
        tck3            : in     vl_logic;
        rlol3           : in     vl_logic;
        rlos_hi3        : in     vl_logic;
        rlos_lo3        : in     vl_logic;
        pci_connect3    : in     vl_logic;
        pci_det_done3   : in     vl_logic;
        refck2core      : in     vl_logic;
        rxrefck2core    : in     vl_logic;
        plol            : in     vl_logic;
        refloc          : in     vl_logic;
        rrefloc         : in     vl_logic;
        rx_ch           : in     vl_logic_vector(3 downto 0);
        scan_out_tx0    : in     vl_logic;
        scan_out_tx1    : in     vl_logic;
        scan_out_tx2    : in     vl_logic;
        scan_out_tx3    : in     vl_logic;
        scan_out_rx0    : in     vl_logic;
        scan_out_rx1    : in     vl_logic;
        scan_out_rx2    : in     vl_logic;
        scan_out_rx3    : in     vl_logic;
        mpif_rd_out     : in     vl_logic_vector(7 downto 0);
        scan_mpif_char_out_prev: in     vl_logic_vector(21 downto 0);
        quad_id         : in     vl_logic_vector(1 downto 0);
        testclk_maco    : in     vl_logic;
        bist_rssigso    : in     vl_logic;
        ubs_bistcomplete: in     vl_logic;
        bist_char_out_prev: in     vl_logic_vector(21 downto 0);
        sds_test_bus    : in     vl_logic_vector(7 downto 0);
        bist_flag_local : in     vl_logic_vector(11 downto 0)
    );
end char_test_logic;
