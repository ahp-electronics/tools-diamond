library verilog;
use verilog.vl_types.all;
entity sram_exec is
    generic(
        AID_SIZE        : integer := 9;
        EA_AUTO         : integer := 10;
        a_width         : integer := 14;
        b_width         : integer := 5;
        DIV             : integer := 29
    );
    port(
        pe_rdata        : out    vl_logic_vector(71 downto 0);
        busy_sram       : out    vl_logic;
        fail_sram       : out    vl_logic;
        sf_be_success   : out    vl_logic;
        sf_ppt_addr     : out    vl_logic_vector(3 downto 0);
        cfg_addr_slew   : out    vl_logic;
        cfg_data_cap    : out    vl_logic;
        cfg_data_flt    : out    vl_logic;
        cfg_data_pre    : out    vl_logic;
        sf_dsr_rst      : out    vl_logic;
        sf_dsr_cap      : out    vl_logic;
        sf_dsr_upd_lat  : out    vl_logic;
        sf_asr_in       : out    vl_logic;
        sf_asr_rst      : out    vl_logic;
        sf_asr_en_incr  : out    vl_logic;
        sf_asr_shift_1st: out    vl_logic;
        sf_asr_shift_2nd: out    vl_logic;
        sf_asr_shift_3rd: out    vl_logic;
        sf_wl_str       : out    vl_logic;
        sf_data_wr      : out    vl_logic;
        sf_es_o         : out    vl_logic_vector(35 downto 0);
        sf_pcs_o        : out    vl_logic_vector(27 downto 0);
        sf_finish_bke   : out    vl_logic;
        jtag_active_smsync: in     vl_logic;
        mc1_bl_float    : in     vl_logic;
        mc1_wl_slew     : in     vl_logic;
        ASR_LENGTH      : in     vl_logic_vector(13 downto 0);
        lsc_done        : in     vl_logic;
        done_gwe        : in     vl_logic;
        lsc_done_ebr    : in     vl_logic;
        lsc_done_ip     : in     vl_logic;
        ctrl_ebr_init_en: in     vl_logic;
        mx_smclk        : in     vl_logic;
        sf_rst_async    : in     vl_logic;
        smclk           : in     vl_logic;
        sf_rst_sync     : in     vl_logic;
        isc_exec_a      : in     vl_logic;
        isc_exec_b      : in     vl_logic;
        isc_exec_c      : in     vl_logic;
        isc_exec_d      : in     vl_logic;
        isc_exec_e      : in     vl_logic;
        isc_exec_f      : in     vl_logic;
        buf128_dat      : in     vl_logic_vector(127 downto 0);
        njpcs_addr_dat  : in     vl_logic_vector(14 downto 0);
        start_bke       : in     vl_logic;
        ebr_init_en     : in     vl_logic;
        sf_prog_exec    : in     vl_logic;
        sf_read_exec    : in     vl_logic;
        sf_erase_exec   : in     vl_logic;
        sf_prog_incr_exec: in     vl_logic;
        sf_read_incr_exec: in     vl_logic;
        sf_pcs_write_exec: in     vl_logic;
        sf_ebr_write_exec: in     vl_logic;
        sf_pcs_read_exec: in     vl_logic;
        sf_ebr_read_exec: in     vl_logic;
        sdm_init_sram_asr_exec: in     vl_logic;
        ppt_init_tsf_asr_exec: in     vl_logic;
        ppt_write_incr_exec: in     vl_logic;
        sf_write_bus_addr_exec: in     vl_logic;
        sf_init_addr_exec: in     vl_logic;
        sf_write_addr_exec: in     vl_logic;
        sf_address_shift_exec: in     vl_logic;
        sed_init_addr_exec: in     vl_logic;
        sed_read_incr_exec: in     vl_logic;
        es_i            : in     vl_logic_vector(8 downto 0);
        pcs_i           : in     vl_logic_vector(7 downto 0);
        pcs_stat        : in     vl_logic_vector(2 downto 0)
    );
end sram_exec;
