library verilog;
use verilog.vl_types.all;
entity regfile is
    port(
        CHIPID          : in     vl_logic_vector(7 downto 0);
        HCLK            : in     vl_logic;
        HRESETn         : in     vl_logic;
        HGRANT_CFG      : in     vl_logic;
        HADDR           : in     vl_logic_vector(17 downto 0);
        HTRANS          : in     vl_logic_vector(1 downto 0);
        HWRITE          : in     vl_logic;
        HSIZE           : in     vl_logic_vector(1 downto 0);
        HWDATAin        : in     vl_logic_vector(31 downto 0);
        HSELExtMem      : in     vl_logic;
        HREADYin        : in     vl_logic;
        HMASTER         : in     vl_logic_vector(3 downto 0);
        RST_LOCK        : in     vl_logic;
        RDATA_READY     : in     vl_logic;
        WDATA_ACK       : in     vl_logic;
        CFG_IRQ_DATA    : in     vl_logic;
        FPSC_BIT_ERR    : in     vl_logic;
        RAM_BIT_ERR     : in     vl_logic;
        ERR_FLAG        : in     vl_logic_vector(1 downto 0);
        RDATA           : in     vl_logic_vector(31 downto 0);
        USER_IRQ_GENERAL: in     vl_logic;
        USER_IRQ_SLAVE  : in     vl_logic;
        USER_IRQ_MASTER : in     vl_logic;
        MPI_IRQ         : in     vl_logic;
        FPSC_IRQ_SLAVE  : in     vl_logic;
        FPSC_IRQ_MASTER : in     vl_logic;
        DEVICE_ID       : in     vl_logic_vector(31 downto 0);
        INTERRUPT_VECTOR_1: in     vl_logic_vector(31 downto 0);
        INTERRUPT_VECTOR_2: in     vl_logic_vector(31 downto 0);
        INTERRUPT_VECTOR_3: in     vl_logic_vector(31 downto 0);
        INTERRUPT_VECTOR_4: in     vl_logic_vector(31 downto 0);
        INTERRUPT_VECTOR_5: in     vl_logic_vector(31 downto 0);
        INTERRUPT_VECTOR_6: in     vl_logic_vector(31 downto 0);
        RDBK_ADDR_ERR   : in     vl_logic;
        CFG_BUS_ERR     : in     vl_logic_vector(1 downto 0);
        BUS_ERR_ADDR    : in     vl_logic_vector(17 downto 0);
        Reset_CFG       : in     vl_logic;
        MC1_MPI         : in     vl_logic;
        MC1_USER        : in     vl_logic;
        MC1_FPSC        : in     vl_logic;
        SCANEN          : in     vl_logic;
        Done            : in     vl_logic;
        InitN           : in     vl_logic;
        MC1_ParityOdd   : in     vl_logic;
        BUS_DATA_LOST   : in     vl_logic;
        BUS_TRAP_ADDR   : in     vl_logic_vector(17 downto 0);
        HRDATAout       : out    vl_logic_vector(35 downto 0);
        HREADYout       : out    vl_logic;
        HRESP           : out    vl_logic_vector(1 downto 0);
        MPI_PAR_CHK     : out    vl_logic;
        PCS_SL_STRAIT   : out    vl_logic;
        MPI_DMA_ENABLE  : out    vl_logic;
        MPI_USR_ENABLE  : out    vl_logic;
        SYS_RD_CFG      : out    vl_logic;
        SYS_GSR         : out    vl_logic;
        PRGM_MPI        : out    vl_logic;
        PRGM_FPSC       : out    vl_logic;
        PRGM_USER       : out    vl_logic;
        SYS_DAISY       : out    vl_logic;
        RDATA_ACK       : out    vl_logic;
        RDATA_SIZE      : out    vl_logic_vector(1 downto 0);
        WDATA_READY     : out    vl_logic;
        WDATA_SIZE      : out    vl_logic_vector(1 downto 0);
        WDATA           : out    vl_logic_vector(31 downto 0);
        RDBK_ADDR       : out    vl_logic_vector(13 downto 0);
        HRESETn_OUT     : out    vl_logic;
        LOCK_FPSC       : out    vl_logic;
        LOCK_USER       : out    vl_logic;
        LOCK_MPI        : out    vl_logic;
        MPI_IRQ_MASKED  : out    vl_logic;
        USER_IRQ_MASKED : out    vl_logic;
        FPSC_IRQ_MASKED : out    vl_logic;
        RFR_EXP         : out    vl_logic_vector(3 downto 0);
        SRI_CLK         : out    vl_logic;
        SRI_RD          : out    vl_logic;
        SRI_WR          : out    vl_logic;
        SRI_RDATA       : in     vl_logic_vector(63 downto 0);
        SRI_WDATA       : out    vl_logic;
        SRI_ADDR        : out    vl_logic_vector(9 downto 0);
        REPEAT_RDBK     : out    vl_logic
    );
end regfile;
