library verilog;
use verilog.vl_types.all;
entity config_inst_dec is
    port(
        instruction     : in     vl_logic_vector(7 downto 0);
        jtag_functional : in     vl_logic;
        edit_mod        : in     vl_logic;
        ee_mod          : in     vl_logic;
        xsram           : in     vl_logic;
        xee             : in     vl_logic;
        edsram          : in     vl_logic;
        edee            : in     vl_logic;
        mfgen           : in     vl_logic;
        rti             : in     vl_logic;
        jtag_unprogram  : in     vl_logic;
        toe             : in     vl_logic;
        mfg_jtag_store  : in     vl_logic;
        mfg_era_red_sel : in     vl_logic;
        mfg_prg_red_sel : in     vl_logic;
        mfg_prg_trim_sel: in     vl_logic;
        goe_high_r      : in     vl_logic;
        tck             : in     vl_logic;
        por             : in     vl_logic;
        mc1_goe_en      : in     vl_logic;
        usr_goe         : in     vl_logic;
        tlreset         : in     vl_logic;
        decrypt_en      : in     vl_logic;
        seldr           : in     vl_logic;
        post_edit       : in     vl_logic;
        done_reg        : in     vl_logic;
        progdis_o       : out    vl_logic;
        progen_ee_o     : out    vl_logic;
        progen_sram_o   : out    vl_logic;
        xprogen_ee_o    : out    vl_logic;
        xreaden_sram_o  : out    vl_logic;
        rst_addr_o      : out    vl_logic;
        erase_ee_o      : out    vl_logic;
        erase_sram_o    : out    vl_logic;
        eraseall_ee_o   : out    vl_logic;
        eraseall_sram_o : out    vl_logic;
        read_o          : out    vl_logic;
        vfy_incr_rti_o  : out    vl_logic;
        ucode_o         : out    vl_logic;
        ucode_ee_o      : out    vl_logic;
        idcode_o        : out    vl_logic;
        selbyp_b        : out    vl_logic;
        selbsr          : out    vl_logic;
        selasr          : out    vl_logic;
        seldsr          : out    vl_logic;
        bsmode1         : out    vl_logic;
        bsmode2         : out    vl_logic;
        bsmode3         : out    vl_logic;
        seler1          : out    vl_logic;
        seler2          : out    vl_logic;
        selid           : out    vl_logic;
        extest          : out    vl_logic;
        sample          : out    vl_logic;
        mnfgshift       : out    vl_logic;
        progee_status   : out    vl_logic;
        readee_status   : out    vl_logic;
        program_ee_o    : out    vl_logic;
        program_sram_o  : out    vl_logic;
        prog_inc_rti_ee_o: out    vl_logic;
        prog_inc_rti_sram_o: out    vl_logic;
        progucode_ee_o  : out    vl_logic;
        progucode_sram_o: out    vl_logic;
        progpes_ee_o    : out    vl_logic;
        progsec_ee_o    : out    vl_logic;
        progsec_sram_o  : out    vl_logic;
        progdone_ee_o   : out    vl_logic;
        progdone_sram_o : out    vl_logic;
        read_pes_o      : out    vl_logic;
        read_ee_o       : out    vl_logic;
        vfy_incr_rti_ee_o: out    vl_logic;
        progctrl0_o     : out    vl_logic;
        vfyctrl0_o      : out    vl_logic;
        refresh_out     : out    vl_logic;
        j_fl_ep         : out    vl_logic;
        j_fl_ep_only    : out    vl_logic;
        mfg_era_red     : out    vl_logic;
        mfg_prg_red     : out    vl_logic;
        read_dnld_red   : out    vl_logic;
        verify_jtag     : out    vl_logic;
        erase_tag_o     : out    vl_logic;
        prog_tag_o      : out    vl_logic;
        read_tag_o      : out    vl_logic;
        jtag_store      : out    vl_logic;
        program_spi     : out    vl_logic;
        progcrc32_o     : out    vl_logic;
        progcrc32_ee_o  : out    vl_logic;
        read_crc_o      : out    vl_logic;
        read_crc_ee_o   : out    vl_logic;
        decrypt_o       : out    vl_logic;
        prog_encr_ee_o  : out    vl_logic;
        read_encr_ee_o  : out    vl_logic;
        erase_encr_ee_o : out    vl_logic;
        protect_shf_o   : out    vl_logic;
        reset_crc16     : out    vl_logic;
        read_crc16      : out    vl_logic;
        encrypt_pgm_inc : out    vl_logic;
        cap_bp          : out    vl_logic;
        red_latch_rst   : out    vl_logic;
        prog_tag        : out    vl_logic;
        read_tag        : out    vl_logic;
        muxclk_en       : out    vl_logic
    );
end config_inst_dec;
