//***************************************************************
// 8-bit up counters with asynchronous clear, CAI, and CAO.
// XiaoQiu ZHOU
//***************************************************************
module CBU18(Q0, Q1, Q2, Q3, Q4, Q5, Q6, Q7, CAO, CAI, CLK, CD);
  output Q0;
  output Q1;
  output Q2;
  output Q3;
  output Q4;
  output Q5;
  output Q6;
  output Q7;
  output CAO;
  input CAI;
  input CLK;
  input CD;
  reg [7:0] Q_i;

always @(posedge CLK or posedge CD)
begin
  if (CD) 
    Q_i = 8'b00000000;		
  else if (CAI) 
    Q_i = Q_i + 1;
end

assign Q0 = Q_i[0];
assign Q1 = Q_i[1];
assign Q2 = Q_i[2];
assign Q3 = Q_i[3];
assign Q4 = Q_i[4];
assign Q5 = Q_i[5];
assign Q6 = Q_i[6];
assign Q7 = Q_i[7];
assign CAO = CAI && Q_i[0] && Q_i[1] && Q_i[2] && Q_i[3] 
&& Q_i[4] && Q_i[5] && Q_i[6] && Q_i[7];

endmodule

