library verilog;
use verilog.vl_types.all;
entity LP0_UDP is
    -- This module cannot be connected to from
    -- VHDL because it has unnamed ports.
end LP0_UDP;
