library verilog;
use verilog.vl_types.all;
entity config_inst_dec is
    port(
        wakeup          : in     vl_logic;
        clear_memory    : in     vl_logic;
        rti             : in     vl_logic;
        instruction     : in     vl_logic_vector(7 downto 0);
        jtag_unprogram  : in     vl_logic;
        jtag_functional : in     vl_logic;
        edit_mod        : in     vl_logic;
        xread_mod       : in     vl_logic;
        post_edit       : in     vl_logic;
        nonjtag_cfg_r   : in     vl_logic;
        read_back_r     : in     vl_logic;
        preamble        : in     vl_logic;
        isc_inst_tri    : out    vl_logic;
        progen          : out    vl_logic;
        progen_o        : out    vl_logic;
        progdis_o       : out    vl_logic;
        xread_en_o      : out    vl_logic;
        xread_dis_o     : out    vl_logic;
        burst_o         : out    vl_logic;
        rst_addr_o      : out    vl_logic;
        erase_o         : out    vl_logic;
        prog_inc_rti_o  : out    vl_logic;
        vfy_incr_rti_o  : out    vl_logic;
        progucode_o     : out    vl_logic;
        ucode_o         : out    vl_logic;
        progctrl0_o     : out    vl_logic;
        vfyctrl0_o      : out    vl_logic;
        rst_crc_o       : out    vl_logic;
        vfy_crc_o       : out    vl_logic;
        progsec_o       : out    vl_logic;
        progdone_o      : out    vl_logic;
        erasedone_o     : out    vl_logic;
        idcode_o        : out    vl_logic;
        status_o        : out    vl_logic;
        ipa_o           : out    vl_logic;
        ipb_o           : out    vl_logic;
        iptesta_o       : out    vl_logic;
        iptestb_o       : out    vl_logic;
        selbyp_b        : out    vl_logic;
        selbsr          : out    vl_logic;
        selasr          : out    vl_logic;
        seldsr          : out    vl_logic;
        bsmode1         : out    vl_logic;
        bsmode2         : out    vl_logic;
        bsmode3         : out    vl_logic;
        test_inst       : out    vl_logic;
        seler1          : out    vl_logic;
        seler2          : out    vl_logic;
        selid           : out    vl_logic;
        nonjtag_active  : out    vl_logic;
        extest          : out    vl_logic;
        sample          : out    vl_logic;
        edit_xread      : out    vl_logic;
        mnfgshift       : out    vl_logic;
        refresh_out     : out    vl_logic
    );
end config_inst_dec;
