library verilog;
use verilog.vl_types.all;
entity CCLK_TREE is
    port(
        A               : in     vl_logic;
        Z               : out    vl_logic
    );
end CCLK_TREE;
