library verilog;
use verilog.vl_types.all;
entity chif is
    generic(
        creg            : integer := 24;
        sreg            : integer := 25
    );
    port(
        pcs_addro       : out    vl_logic_vector(7 downto 0);
        pcs_rdo         : out    vl_logic;
        pcs_wdatao      : out    vl_logic_vector(7 downto 0);
        pcs_wstbo       : out    vl_logic;
        pcs_rdata_qxcyo : out    vl_logic_vector(7 downto 0);
        pcs_into        : out    vl_logic;
        start_seq_wstr  : out    vl_logic;
        a1a2_mpi_wstr   : out    vl_logic;
        b1_mpi_wstr     : out    vl_logic;
        k2_mpi_wstr     : out    vl_logic;
        set_np_loaded_wstr: out    vl_logic;
        int_cha_out     : out    vl_logic;
        gen_ctl_1_ba_00 : out    vl_logic_vector(7 downto 0);
        gen_ctl_2_ba_01 : out    vl_logic_vector(7 downto 0);
        gen_ctl_3_ba_02 : out    vl_logic_vector(7 downto 0);
        pkt_ctl_1_ba_05 : out    vl_logic_vector(7 downto 0);
        pkt_ctl_2_ba_06 : out    vl_logic_vector(7 downto 0);
        pkt_ctl_3_ba_07 : out    vl_logic_vector(7 downto 0);
        pkt_ctl_4_ba_08 : out    vl_logic_vector(7 downto 0);
        pkt_ctl_5_ba_09 : out    vl_logic_vector(7 downto 0);
        son_ctl_1_ba_0b : out    vl_logic_vector(7 downto 0);
        son_ctl_2_ba_0c : out    vl_logic_vector(7 downto 0);
        son_ctl_3_ba_0d : out    vl_logic_vector(7 downto 0);
        son_ctl_4_ba_0e : out    vl_logic_vector(7 downto 0);
        son_ctl_5_ba_0f : out    vl_logic_vector(7 downto 0);
        son_ctl_6_ba_10 : out    vl_logic_vector(7 downto 0);
        son_ctl_7_ba_11 : out    vl_logic_vector(7 downto 0);
        ser_ctl_1_ba_13 : out    vl_logic_vector(7 downto 0);
        ser_ctl_2_ba_14 : out    vl_logic_vector(7 downto 0);
        ser_ctl_3_ba_15 : out    vl_logic_vector(7 downto 0);
        ser_ctl_4_ba_16 : out    vl_logic_vector(7 downto 0);
        pcs_inti        : in     vl_logic;
        resetn          : in     vl_logic;
        pcs_addri       : in     vl_logic_vector(7 downto 0);
        pcs_wdatai      : in     vl_logic_vector(7 downto 0);
        pcs_wstbi       : in     vl_logic;
        pcs_rdi         : in     vl_logic;
        pcs_qxcyi       : in     vl_logic;
        pcs_rdata_qxcyi : in     vl_logic_vector(7 downto 0);
        test_clk        : in     vl_logic;
        test_mode       : in     vl_logic;
        force_int       : in     vl_logic;
        prbs_error      : in     vl_logic;
        bip_error       : in     vl_logic;
        gen_sts_1_ba_80 : in     vl_logic_vector(7 downto 0);
        gen_sts_3_ba_82 : in     vl_logic_vector(7 downto 0);
        gen_sts_4_ba_83 : in     vl_logic_vector(7 downto 0);
        pkt_sts_1_ba_85 : in     vl_logic_vector(7 downto 0);
        pkt_sts_2_ba_86 : in     vl_logic_vector(7 downto 0);
        pkt_sts_3_ba_87 : in     vl_logic_vector(7 downto 0);
        pkt_sts_4_ba_88 : in     vl_logic_vector(7 downto 0);
        pkt_sts_5_ba_89 : in     vl_logic_vector(7 downto 0);
        son_sts_1_ba_8b : in     vl_logic_vector(7 downto 0);
        son_sts_3_ba_8d : in     vl_logic_vector(7 downto 0);
        son_sts_4_ba_8e : in     vl_logic_vector(7 downto 0);
        son_sts_5_ba_8f : in     vl_logic_vector(7 downto 0);
        son_sts_6_ba_90 : in     vl_logic_vector(7 downto 0);
        son_sts_7_ba_91 : in     vl_logic_vector(7 downto 0);
        son_sts_8_ba_92 : in     vl_logic_vector(7 downto 0);
        ser_sts_1_ba_94 : in     vl_logic_vector(7 downto 0);
        ser_sts_2_ba_95 : in     vl_logic_vector(7 downto 0);
        ser_sts_3_ba_96 : in     vl_logic_vector(7 downto 0)
    );
end chif;
