module ICC(
TXCLK, TXREADY, TXVALID, TXDATA0, TXDATA1, TXDATA2,
TXDATA3, TXDATA4, TXDATA5, TXDATA6, TXDATA7, INT,
AUX, TXVIO0, TXVIO1, RXVIO0, RXVIO1, RXCLK, RXREADY,
RXVALID, RXDATA0, RXDATA1, RXDATA2, RXDATA3, RXDATA4,
RXDATA5, RXDATA6, RXDATA7);

input TXCLK, TXREADY, TXVALID, TXDATA0, TXDATA1, TXDATA2;
input TXDATA3, TXDATA4, TXDATA5, TXDATA6, TXDATA7, INT;
input AUX, TXVIO0, TXVIO1;

output RXVIO0, RXVIO1, RXCLK, RXREADY;
output RXVALID, RXDATA0, RXDATA1, RXDATA2, RXDATA3, RXDATA4;
output RXDATA5, RXDATA6, RXDATA7;


assign RXVIO0	=	1'b0;
assign RXVIO1   =	1'b0;
assign RXCLK    =	1'b0;
assign RXREADY  =	1'b0;
assign RXVALID  =	1'b0;
assign RXDATA0  =	1'b0;
assign RXDATA1  =	1'b0;
assign RXDATA2  =	1'b0;
assign RXDATA3  =	1'b0;
assign RXDATA4  =	1'b0;
assign RXDATA5  =	1'b0;
assign RXDATA6  =	1'b0;
assign RXDATA7  =	1'b0;

endmodule