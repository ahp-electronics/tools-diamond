library verilog;
use verilog.vl_types.all;
entity SSPIA is
    generic(
        TAG_INITSIZE    : integer := 2184;
        TAG_INITVAL_00  : string  := "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
        TAG_INITVAL_01  : string  := "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
        TAG_INITVAL_02  : string  := "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
        TAG_INITVAL_03  : string  := "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
        TAG_INITVAL_04  : string  := "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
        TAG_INITVAL_05  : string  := "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
        TAG_INITVAL_06  : string  := "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
        TAG_INITVAL_07  : string  := "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
        TAG_INITVAL_08  : string  := "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
        TAG_INITVAL_09  : string  := "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
        TAG_INITVAL_0A  : string  := "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
        TAG_INITVAL_0B  : string  := "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
        TAG_INITVAL_0C  : string  := "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000"
    );
    port(
        SI              : in     vl_logic;
        CLK             : in     vl_logic;
        CS              : in     vl_logic;
        SO              : out    vl_logic
    );
end SSPIA;
