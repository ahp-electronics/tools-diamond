--
@ER--B$FbsEHo0OR52gR4g-cRRj.jd$R1MHbDO$H0ROQM
R--fN]C8:CsR#//$DMbH0OH$N/lb..jjDjdNl0/NCbbsG#/HMDHGH/DLC/oMHCsOC/oMC_oMHCsON/slI_sb3_sPyE84
Rf-
-
----- RBpXpR)dqv.7X4R----D-
HNLssH$RC;CC
Ck#RCHCC03#8F_Do_HO4c4n3DND;#
kCCRHC#C30D8_FOoH_o#HM3C8N;DD
LDHs$NsRHkM#;Hl
Ck#RHkM#3HlPlOFbCFMM30#N;DD
M
C0$H0RqX)vXd.4H7R#R
Rb0FsRR5
RRRRR7RRuRmRRF:Rk#0R0k8_DHFoOR;RRRRRRRR
RRRRR1RRuRmRRF:Rk#0R0k8_DHFoO
;
RRRRRRRRqRjRRRR:H#MR0k8_DHFoOR;
RRRRRqRR4RRRRH:RM0R#8D_kFOoH;R
RRRRRR.RqRRRR:MRHR8#0_FkDo;HO
RRRRRRRRRqdR:RRRRHM#_08koDFH
O;RRRRRRRRqRcRRRR:H#MR0k8_DHFoOR;
RRRRR7RRRRRRRH:RM0R#8D_kFOoH;R
RRRRRRuR7)Rqj:MRHR8#0_FkDo;HO
RRRRRRRR)7uq:4RRRHM#_08koDFH
O;RRRRRRRR7qu).RR:H#MR0k8_DHFoOR;
RRRRR7RRud)qRH:RM0R#8D_kFOoH;R
RRRRRRuR7)Rqc:MRHR8#0_FkDo;HO
RRRRRRRRpWBi:RRRRHM#_08koDFHRO;RRRRR
RRRRRRRRRRWR RRRR:H#MR0k8_DHFoOR
RRRRRRR2;RM
C8)RXq.vdX;47
ONsECH0Os0kC)RXq.vdX_47eVRFRqX)vXd.4H7R#R
RSo#HMRNDI,CjR4IC,FR#j#,RFR4,8,FjR48F:0R#8F_Do;HO
oLCHSM
7Rum<8=RFIjRERCM5)7uq=cRR''j2DRC#8CRF
4;Sm1uRR<=#RFjIMECRc5qR'=RjR'2CCD#R4#F;I
SC<jR= RWR8NMRF5M0cRq2S;
IRC4<W=R MRN8cRq;S
Rz:jRRv)q44nX7RR
RRRRRRRRRRRRRbRRFRs0lRNb5=7R>,R7RRqj=q>Rjq,R4>R=R,q4RRq.=q>R.q,Rd>R=R,qd
SRSS)7uq=jR>uR7),qjR)7uq=4R>uR7),q4R)7uq=.R>uR7),q.R)7uq=dR>uR7),qdRS
SSRW =I>RCRj,WiBpRR=>WiBp,uR7m>R=Rj8F,uR1m>R=Rj#F2R;
SRz4:qR)vX4n4
7RRRRRRRRRRRRRRRRRb0FsRblNRR57=7>R,jRqRR=>qRj,q=4R>4Rq,.RqRR=>qR.,q=dR>dRq,S
RSuS7)Rqj=7>Ruj)q,uR7)Rq4=7>Ru4)q,uR7)Rq.=7>Ru.)q,uR7)Rqd=7>Rud)q,SR
S SWRR=>I,C4RpWBi>R=RpWBi7,Ru=mR>FR841,Ru=mR>FR#4
2;CRM8Xv)qd4.X7;_e
-
--R--Bp pRqX)vXnc4-7R----
LDHs$NsRCHCCk;
#HCRC3CC#_08DHFoO4_4nNc3D
D;kR#CHCCC38#0_oDFH#O_HCoM8D3NDD;
HNLssk$RMHH#lk;
#kCRMHH#lO3PFFlbM0CM#D3ND
;
CHM00X$R)nqvc7X4R
H#RFRbs50R
RRRRRRRRm7uR:RRR0FkR8#0_FkDo;HORRRRRRRR
RRRRRRRRm1uR:RRR0FkR8#0_FkDo;HO
R
RRRRRRjRqRRRR:MRHR8#0_FkDo;HO
RRRRRRRRRq4R:RRRRHM#_08koDFH
O;RRRRRRRRqR.RRRR:H#MR0k8_DHFoOR;
RRRRRqRRdRRRRH:RM0R#8D_kFOoH;R
RRRRRRcRqRRRR:MRHR8#0_FkDo;HO
RRRRRRRRRq6R:RRRRHM#_08koDFH
O;RRRRRRRR7RRRRRR:H#MR0k8_DHFoOR;
RRRRR7RRuj)qRH:RM0R#8D_kFOoH;R
RRRRRRuR7)Rq4:MRHR8#0_FkDo;HO
RRRRRRRR)7uq:.RRRHM#_08koDFH
O;RRRRRRRR7qu)dRR:H#MR0k8_DHFoOR;
RRRRR7RRuc)qRH:RM0R#8D_kFOoH;R
RRRRRRuR7)Rq6:MRHR8#0_FkDo;HO
RRRRRRRRpWBi:RRRRHM#_08koDFHRO;RRRRR
RRRRRRRRRRWR RRRR:H#MR0k8_DHFoOR
RRRRRRR2;RM
C8)RXqcvnX;47
ONsECH0Os0kC)RXqcvnX_47eVRFRqX)vXnc4H7R#R
RSo#HMRNDI,CjR4IC,CRI.I,RCRd,#,FjR4#F,FR#.#,RFRd,8,FjR48F,FR8.8,RFRd:#_08DHFoOL;
CMoH
uS7m=R<RFR8jERIC5MR7qu)6RR='Rj'NRM87qu)cRR='2j'R#CDCSR
S48FRCIEM7R5u6)qR'=RjN'RM78Ruc)qR'=R4R'2CCD#RS
S8RF.IMECRu57)Rq6=4R''MRN8uR7)Rqc=jR''C2RDR#C
8SSF
d;Sm1uRR<=Rj#FRCIEMqR56RR='Rj'NRM8q=cRR''j2DRC#
CRSFS#4ERIC5MRq=6RR''jR8NMRRqc=4R''C2RDR#C
#SSFI.RERCM5Rq6=4R''MRN8cRqR'=RjR'2CCD#RS
S#;Fd
CSIj=R<RRW NRM850MFR2q6R8NMRF5M0cRq2S;
IRC4<W=R MRN8MR5Fq0R6N2RMq8RcS;
IRC.<W=R MRN86RqR8NMRF5M0cRq2S;
IRCd<W=R MRN86RqR8NMR;qc
zRSjRR:)4qvn7X4RR
RRRRRRRRRRRRRRFRbsl0RN5bR7>R=RR7,q=jR>jRq,4RqRR=>qR4,q=.R>.Rq,dRqRR=>q
d,RSSS7qu)j>R=R)7uqRj,7qu)4>R=R)7uqR4,7qu).>R=R)7uqR.,7qu)d>R=R)7uqRd,
SSSW= R>CRIjW,RBRpi=W>RB,piRm7uRR=>8,FjRm1uRR=>#2Fj;S
Rz:4RRv)q44nX7RR
RRRRRRRRRRRRRbRRFRs0lRNb5=7R>,R7RRqj=q>Rjq,R4>R=R,q4RRq.=q>R.q,Rd>R=R,qd
SRSS)7uq=jR>uR7),qjR)7uq=4R>uR7),q4R)7uq=.R>uR7),q.R)7uq=dR>uR7),qdRS
SSRW =I>RCR4,WiBpRR=>WiBp,uR7m>R=R48F,uR1m>R=R4#F2R;
SRz.:qR)vX4n4
7RRRRRRRRRRRRRRRRRb0FsRblNRR57=7>R,jRqRR=>qRj,q=4R>4Rq,.RqRR=>qR.,q=dR>dRq,S
RSuS7)Rqj=7>Ruj)q,uR7)Rq4=7>Ru4)q,uR7)Rq.=7>Ru.)q,uR7)Rqd=7>Rud)q,SR
S SWRR=>I,C.RpWBi>R=RpWBi7,Ru=mR>FR8.1,Ru=mR>FR#.
2;RdSzR):Rqnv4XR47
RRRRRRRRRRRRRRRRsbF0NRlb7R5RR=>7q,Rj>R=R,qjRRq4=q>R4q,R.>R=R,q.RRqd=q>RdR,
S7SSuj)qRR=>7qu)j7,Ru4)qRR=>7qu)47,Ru.)qRR=>7qu).7,Rud)qRR=>7qu)d
,RSWSS >R=RdIC,BRWp=iR>BRWpRi,7Rum=8>RFRd,1Rum=#>RF;d2
8CMRqX)vXnc4e7_;-

--
-
R--1bHlD)CRqIvRHR0E#oHMDqCR7 7)1V1RFLsRFR0Es8CNR8NMRHIs0-C
-NRas0oCRX:RHMDHG-
-
H
DLssN$CRHC
C;kR#CHCCC38#0_oDFH4O_43ncN;DD
Ck#RCHCC03#8F_Do_HO#MHoCN83D
D;DsHLNRs$k#MHH
l;kR#Ck#MHHPl3ObFlFMMC0N#3D
D;CHM00)$Rq)v_W)u_R
H#SMoCCOsHRS5
RRRRVHNlD:$RRs#0HRMo:"=RMCFM"S;
S8IH0:ERR0HMCsoCRR:=4
;RS8SN8HsI8R0E:MRH0CCos=R:RRn;RRRRR-RR-HRLoMRCFEkoRsVFRb8C0SE
Sb8C0:ERR0HMCsoCRR:=c
U;S8SsF_k0sRCo:FRLFNDCM=R:RDVN#RC;RRRRRR--ERN#Fbk0ks0RCSo
SFI8ks0_C:oRRFLFDMCNRR:=V#NDCS;S-E-RNF#Rkk0b0CRsoS
S8_HMsRCo:FRLFNDCM=R:RDVN#RC;RRRRR-RR-NRE#NR80HNRM0bkRosC
sSSNs88_osCRL:RFCFDN:MR=NRVD;#CRRRRR-R-R#ENRNsC88RN8#sC#CRsoS
SI8N8sC_soRR:LDFFCRNMRR:=V#NDCRRRR-RR-NRE#sRIHR0CNs88CR##s
CoS;S2
FSbs50R
)SS_z7maF:Rk#0R0D8_FOoH_OPC05FsI0H8ER-48MFI0jFR2S;
S7W_mRza:kRF00R#8F_Do_HOP0COFIs5HE80-84RF0IMF2Rj;S
S)7q7)RR:H#MR0D8_FOoH_OPC05FsNs88I0H8ER-48MFI0jFR2S;
Sh7QRRR:H#MR0D8_FOoH_OPC05FsI0H8ER-48MFI0jFR2S;
S7Wq7:)RRRHM#_08DHFoOC_POs0F58N8s8IH04E-RI8FMR0Fj
2;S SWRRR:H#MR0D8_FOoH;RRRRRRR-I-RsCH0RNCMLRDCVRFss
NlSpSBiRR:H#MR0D8_FOoH;RRRRRRR-O-RD	FORsVFRlsN,8RN8Rs,8
HMS_S)miBpRH:RM0R#8F_Do;HORRRRR-RR-bRF0DROFRO	VRFssF_8kS0
SmW_BRpi:MRHR8#0_oDFHROR-b-F0FRVs_RI80Fk
2SS;M
C8MRC0$H0Rv)q_u)W_
);

---w-RH0s#RbHlDCClM00NHRFMl0k#RRLCODNDCN8RsjOE

--NEsOHO0C0CksRFLDOs	_NFlRVqR)vW_)uR_)HO#
FFlbM0CMRqX)vXd.4R7RRsbF0
R5RRRRRRRR7RumRRR:FRk0#_08koDFHRO;RRRRR
RRRRRRRRRR1RumRRR:FRk0#_08koDFH
O;
RRRRRRRRRqjR:RRRRHM#_08koDFH
O;RRRRRRRRqR4RRRR:H#MR0k8_DHFoOR;
RRRRRqRR.RRRRH:RM0R#8D_kFOoH;R
RRRRRRdRqRRRR:MRHR8#0_FkDo;HO
RRRRRRRRRqcR:RRRRHM#_08koDFH
O;RRRRRRRR7RRRRRR:H#MR0k8_DHFoOR;
RRRRR7RRuj)qRH:RM0R#8D_kFOoH;R
RRRRRRuR7)Rq4:MRHR8#0_FkDo;HO
RRRRRRRR)7uq:.RRRHM#_08koDFH
O;RRRRRRRR7qu)dRR:H#MR0k8_DHFoOR;
RRRRR7RRuc)qRH:RM0R#8D_kFOoH;R
RRRRRRBRWpRiR:MRHR8#0_FkDo;HORRRRRRRR
RRRRRRRRRW R:RRRRHM#_08koDFHRO
RRRRR;R2RCR
MO8RFFlbM0CM;F
OlMbFCRM0Xv)qn4cX7RRRb0FsRR5
RRRRR7RRuRmRRF:Rk#0R0k8_DHFoOR;RRRRRRRR
RRRRR1RRuRmRRF:Rk#0R0k8_DHFoO
;
RRRRRRRRqRjRRRR:H#MR0k8_DHFoOR;
RRRRRqRR4RRRRH:RM0R#8D_kFOoH;R
RRRRRR.RqRRRR:MRHR8#0_FkDo;HO
RRRRRRRRRqdR:RRRRHM#_08koDFH
O;RRRRRRRRqRcRRRR:H#MR0k8_DHFoOR;
RRRRRqRR6RRRRH:RM0R#8D_kFOoH;R
RRRRRRRR7RRRR:MRHR8#0_FkDo;HO
RRRRRRRR)7uq:jRRRHM#_08koDFH
O;RRRRRRRR7qu)4RR:H#MR0k8_DHFoOR;
RRRRR7RRu.)qRH:RM0R#8D_kFOoH;R
RRRRRRuR7)Rqd:MRHR8#0_FkDo;HO
RRRRRRRR)7uq:cRRRHM#_08koDFH
O;RRRRRRRR7qu)6RR:H#MR0k8_DHFoOR;
RRRRRWRRBRpiRH:RM0R#8D_kFOoH;RRRRRRRRR
RRRRRR RWRRRR:MRHR8#0_FkDo
HORRRRR2RR;
RRCRM8ObFlFMMC0V;
k0MOHRFMVOkM_HHM0R5L:FRLFNDCMs2RCs0kM0R#soHMR
H#LHCoMR
RH5VRL02RE
CMRRRRskC0s"M5"
2;RDRC#RC
RsRRCs0kMB5"F8kDR0MFRbHlDCClMA0RD	FORv)q3#RQRC0ERNsC88RN8#sC#CRso0H#C8sCRHk#M0oRE#CRNRlCOODF	#RNRC0ERv)q?;"2
CRRMH8RVC;
MV8Rk_MOH0MH;k
VMHO0FoMRCC0_M88_CEb05x#HCRR:HCM0oRCs;CR8bR0E:MRH0CCoss2RCs0kMMRH0CCos#RH
sPNHDNLCHRlMH_#x:CRR0HMCsoCRR:=jL;
CMoH
lRRH#M_HRxC:8=RCEb0;R
RH5VR#CHxR8<RCEb02ER0CRM
RlRRH#M_HRxC:#=RH;xC
CRRMH8RVR;
R0sCkRsMl_HM#CHx;M
C8CRo0M_C8C_8b;0E
0N0skHL0oCRCsMCNs0F_bsCFRs0:0R#soHM;0
N0LsHkR0CoCCMsFN0sC_sb0FsRRFVLODF	N_slRR:NEsOHO0C0CksRRH#VOkM_HHM0N5s8_8ss2Co;-
-RoLCHLMRD	FORlsNRbHlDCClM00NHRFM#MHoN
D#0C$bR0HM_sNsNH$R#sRNsRN$50jRF2R6RRFVHCM0o;Cs
MOF#M0N0HRI8_0ENNss$RR:H_M0NNss$=R:R,54RR.,cg,R,UR4,nRd2O;
F0M#NRM080CbEs_NsRN$:MRH0s_NsRN$:5=R4UndcU,R4,g.Rgcjn.,Rj,cUR.4jc6,R4;.2
MOF#M0N0HR8PRd.:MRH0CCos=R:RH5I8-0E4d2/nO;
F0M#NRM084HPnRR:HCM0oRCs:5=RI0H8E2-4/;4U
MOF#M0N0HR8P:URR0HMCsoCRR:=58IH04E-2;/g
MOF#M0N0HR8P:cRR0HMCsoCRR:=58IH04E-2;/c
MOF#M0N0HR8P:.RR0HMCsoCRR:=58IH04E-2;/.
MOF#M0N0HR8P:4RR0HMCsoCRR:=58IH04E-2;/4
F
OMN#0ML0RF4FDRL:RFCFDN:MR=8R5HRP4>2Rj;F
OMN#0ML0RF.FDRL:RFCFDN:MR=8R5HRP.>2Rj;F
OMN#0ML0RFcFDRL:RFCFDN:MR=8R5HRPc>2Rj;F
OMN#0ML0RFUFDRL:RFCFDN:MR=8R5HRPU>2Rj;F
OMN#0ML0RF4FDnRR:LDFFCRNM:5=R84HPnRR>j
2;O#FM00NMRFLFDRd.:FRLFNDCM=R:RH58PRd.>2Rj;O

F0M#NRM084HPncdURH:RMo0CC:sR=8R5CEb0-/424UndcO;
F0M#NRM08UHP4Rg.:MRH0CCos=R:RC58b-0E4U2/4;g.
MOF#M0N0HR8PgcjnRR:HCM0oRCs:5=R80CbE2-4/gcjnO;
F0M#NRM08.HPjRcU:MRH0CCos=R:RC58b-0E4.2/j;cU
MOF#M0N0HR8P.4jcRR:HCM0oRCs:5=R80CbE2-4/.4jcO;
F0M#NRM086HP4:.RR0HMCsoCRR:=5b8C04E-24/6.
;
O#FM00NMRFLFD.64RL:RFCFDN:MR=8R5H4P6.RR>j
2;O#FM00NMRFLFD.4jcRR:LDFFCRNM:5=R84HPjR.c>2Rj;F
OMN#0ML0RF.FDjRcU:FRLFNDCM=R:RH58Pc.jURR>j
2;O#FM00NMRFLFDgcjnRR:LDFFCRNM:5=R8cHPjRgn>2Rj;F
OMN#0ML0RFUFD4Rg.:FRLFNDCM=R:RH58PgU4.RR>j
2;O#FM00NMRFLFDd4nU:cRRFLFDMCNRR:=5P8H4UndcRR>j
2;
MOF#M0N0kR#lH_I8R0E:MRH0CCos=R:RmAmph q'#bF5FLFDR42+mRAmqp hF'b#F5LF2D.RA+Rm mpqbh'FL#5FcFD2RR+Apmm 'qhb5F#LDFFU+2RRmAmph q'#bF5FLFD24n;F
OMN#0M#0Rk8l_CEb0RH:RMo0CC:sR=RR6-AR5m mpqbh'FL#5F6FD4R.2+mRAmqp hF'b#F5LFjD4.Rc2+mRAmqp hF'b#F5LFjD.cRU2+mRAmqp hF'b#F5LFjDcgRn2+mRAmqp hF'b#F5LF4DUg2.2;O

F0M#NRM0IE_OFCHO_8IH0:ERR0HMCsoCRR:=I0H8Es_Ns5N$#_klI0H8E
2;O#FM00NMROI_EOFHCC_8bR0E:MRH0CCos=R:Rb8C0NE_s$sN5l#k_8IH0;E2
MOF#M0N0_R8OHEFOIC_HE80RH:RMo0CC:sR=HRI8_0ENNss$k5#lC_8b20E;F
OMN#0M80R_FOEH_OC80CbERR:HCM0oRCs:8=RCEb0_sNsN#$5k8l_CEb02
;
O#FM00NMRII_HE80_lMk_DOCD:#RR0HMCsoCRR:=58IH04E-2_/IOHEFOIC_HE80R4+R;F
OMN#0MI0R_b8C0ME_kOl_C#DDRH:RMo0CC:sR=8R5CEb0-/42IE_OFCHO_b8C0+ERR
4;
MOF#M0N0_R8I0H8Ek_MlC_ODRD#:MRH0CCos=R:RH5I8-0E482/_FOEH_OCI0H8ERR+4O;
F0M#NRM08C_8b_0EM_klODCD#RR:HCM0oRCs:5=R80CbE2-4/O8_EOFHCC_8bR0E+;R4
F
OMN#0MI0R_x#HCRR:HCM0oRCs:I=R_8IH0ME_kOl_C#DDRI*R_b8C0ME_kOl_C#DD;F
OMN#0M80R_x#HCRR:HCM0oRCs:8=R_8IH0ME_kOl_C#DDR8*R_b8C0ME_kOl_C#DD;O

F0M#NRM0LDFF_:8RRFLFDMCNRR:=5#8_HRxC-_RI#CHxRR<=j
2;O#FM00NMRFLFDR_I:FRLFNDCM=R:R0MF5FLFD2_8;O

F0M#NRM0OHEFOIC_HE80RH:RMo0CC:sR=AR5m mpqbh'FL#5F_FD8*2RRO8_EOFHCH_I820ER5+RApmm 'qhb5F#LDFF_RI2*_RIOHEFOIC_HE802O;
F0M#NRM0OHEFO8C_CEb0RH:RMo0CC:sR=AR5m mpqbh'FL#5F_FD8*2RRO8_EOFHCC_8b20ER5+RApmm 'qhb5F#LDFF_RI2*_RIOHEFO8C_CEb02O;
F0M#NRM0I0H8Ek_MlC_ODRD#:MRH0CCos=R:Rm5Amqp hF'b#F5LF8D_25R*I0H8E2-4/O8_EOFHCH_I820ER5+RApmm 'qhb5F#LDFF_RI2*IR5HE80-/42IE_OFCHO_8IH0RE2+;R4
MOF#M0N0CR8b_0EM_klODCD#RR:HCM0oRCs:5=RApmm 'qhb5F#LDFF_R82*C58b-0E482/_FOEH_OC80CbE+2RRm5Amqp hF'b#F5LFID_2RR*5b8C04E-2_/IOHEFO8C_CEb02RR+40;
$RbCF_k0L4k#_b0$C#RHRsNsN5$R80CbEk_MlC_OD-D#4FR8IFM0RRj,I0H8Ek_MlC_OD-D#4FR8IFM0RRj2F#VR0D8_FOoH;H
#oDMNRksF0k_L#:4RR0Fk_#Lk4$_0bRC;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-7R.RsNsNF$RV_Rs80FkRM5HbRk000FRs#H-0CN0##2
HNoMDFRIkL0_kR#4:kRF0k_L#04_$;bC
b0$CkRF0k_L#0._$RbCHN#Rs$sNRC58b_0EM_klODCD#R-48MFI0jFR,*R.I0H8Ek_MlC_OD+D#4FR8IFM0RRj2F#VR0D8_FOoH;H
#oDMNRksF0k_L#:.RR0Fk_#Lk.$_0bRC;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-7R.RsNsNF$RV_Rs80FkRM5HbRk000FRs#H-0CN0##2
HNoMDFRIkL0_kR#.:kRF0k_L#0._$;bC
b0$CkRF0k_L#0c_$RbCHN#Rs$sNRC58b_0EM_klODCD#R-48MFI0jFR,*RcI0H8Ek_MlC_OD+D#dFR8IFM0RRj2F#VR0D8_FOoH;H
#oDMNRksF0k_L#:cRR0Fk_#Lkc$_0bRC;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-7R.RsNsNF$RV_Rs80FkRM5HbRk000FRs#H-0CN0##2
HNoMDFRIkL0_kR#c:kRF0k_L#0c_$;bC
b0$CkRF0k_L#0U_$RbCHN#Rs$sNRC58b_0EM_klODCD#R-48MFI0jFR,*RUI0H8Ek_MlC_OD+D#(FR8IFM0RRj2F#VR0D8_FOoH;H
#oDMNRksF0k_L#:URR0Fk_#LkU$_0bRC;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-7R.RsNsNF$RV_Rs80FkRM5HbRk000FRs#H-0CN0##2
HNoMDFRIkL0_kR#U:kRF0k_L#0U_$;bC
b0$CNRbs$H0_#LkU$_0bHCR#sRNsRN$5b8C0ME_kOl_C#DD-84RF0IMF,RjR8IH0ME_kOl_C#DD-84RF0IMF2RjRRFV#_08DHFoO#;
HNoMDbRsN0sH$k_L#:URRsbNH_0$LUk#_b0$CR;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-.-R7sRNsRN$FsVR_k8F0HR5M0bkRR0F0-sH#00NC
#2#MHoNIDRbHNs0L$_kR#U:NRbs$H0_#LkU$_0b
C;0C$bR0Fk_#Lk40n_$RbCHN#Rs$sNRC58b_0EM_klODCD#R-48MFI0jFR,nR4*8IH0ME_kOl_C#DD+R468MFI0jFR2VRFR8#0_oDFH
O;#MHoNsDRF_k0L4k#nRR:F_k0L4k#n$_0bRC;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--.N7Rs$sNRRFVsF_8k50RHkMb0FR0RH0s-N#002C#
o#HMRNDI0Fk_#Lk4:nRR0Fk_#Lk40n_$;bC
b0$CNRbs$H0_#Lk40n_$RbCHN#Rs$sNRC58b_0EM_klODCD#R-48MFI0jFR,*R.I0H8Ek_MlC_OD+D#4FR8IFM0RRj2F#VR0D8_FOoH;H
#oDMNRNsbs$H0_#Lk4:nRRsbNH_0$L4k#n$_0bRC;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-7R.RsNsNF$RV_Rs80FkRM5HbRk000FRs#H-0CN0##2
HNoMDbRIN0sH$k_L#R4n:NRbs$H0_#Lk40n_$;bC
b0$CkRF0k_L#_d.0C$bRRH#NNss$8R5CEb0_lMk_DOCD4#-RI8FMR0Fjd,R.H*I8_0EM_klODCD#4+dRI8FMR0FjF2RV0R#8F_Do;HO
o#HMRNDs0Fk_#Lkd:.RR0Fk_#Lkd0._$;bCRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RR.7NNss$VRFR8s_FRk05bHMk00RFsR0H0-#N#0C2H
#oDMNRkIF0k_L#Rd.:kRF0k_L#_d.0C$b;$
0bbCRN0sH$k_L#_d.0C$bRRH#NNss$8R5CEb0_lMk_DOCD4#-RI8FMR0Fjc,R*8IH0ME_kOl_C#DD+8dRF0IMF2RjRRFV#_08DHFoO#;
HNoMDbRsN0sH$k_L#Rd.:NRbs$H0_#Lkd0._$;bCRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-.-R7sRNsRN$FsVR_k8F0HR5M0bkRR0F0-sH#00NC
#2#MHoNIDRbHNs0L$_k.#dRb:RN0sH$k_L#_d.0C$b;H
#oDMNRksF0M_CR#:R0D8_FOoH_OPC05Fs80CbEk_MlC_OD-D#4FR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--CLMNDRC#VRFs0-sH#00NC##
HNoMDFRIkC0_MRR:#_08DHFoOC_POs0F5b8C0ME_kOl_C#DD-84RF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RNCML#DCRsVFRH0s-N#00
C##MHoNIDRsC0_MRR:#_08DHFoOC_POs0F5b8C0ME_kOl_C#DD-84RF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RHIs0CCRMDNLCV#RFCsRNROEsRFIF)VRqOvRC#DD
o#HMRNDHsM_C:oRR8#0_oDFHPO_CFO0sH5I8+0Ed86RF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-k-R#RC80sFRC#oH0RCs7RQh
o#HMRNDs0Fk_osCR#:R0D8_FOoH_OPC05FsI0H8E6+dRI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--k8#CRR0FsHCo#s0CRz7maH
#oDMNRkIF0C_soRR:#_08DHFoOC_POs0F58IH0dE+6FR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RCk#8FR0RosCHC#0smR7z#a
HNoMDFRsks0_CRo4:0R#8F_Do_HOP0COFIs5HE80-84RF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RCk#8FR0RFOEFR#CLIC0CRCM7RQhNRM8Fbk0kF0RVDRAFRO	)
qv#MHoNsDRNs8_C:oRR8#0_oDFHPO_CFO0s85N8HsI8-0E4FR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-#RkC08RFCRso0H#C)sRq)77
o#HMRNDI_N8sRCo:0R#8F_Do_HOP0COFNs58I8sHE80-84RF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-k-R#RC80sFRC#oH0RCsW7q7)H
#oDMNRIDF_8sN8:sRR8#0_oDFHPO_CFO0sd54RI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-R8sN8LsRHR0#HkMb0FR0Rv)qRDOCD5#RcHRL0s#RCHJks2C8
o#HMRNDD_FII8N8sRR:#_08DHFoOC_POs0F5R4d8MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--I8N8sHRL0H#RM0bkRR0F)RqvODCD#cR5R0LH#CRsJskHC
82#MHoN)DRq)77_b0lR#:R0D8_FOoH_OPC05FsNs88I0H8ER-48MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--k8#CRR0FbCHbDCHMR7)q7#)
HNoMDqRW7_7)0Rlb:0R#8F_Do_HOP0COFNs58I8sHE80-84RF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-k-R#RC80bFRHDbCHRMCW7q7)H
#oDMNRh7Q_b0lR#:R0D8_FOoH_OPC05FsI0H8ER-48MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-#RkC08RFHRbbHCDM7CRQ#h
HNoMD RW_b0lR#:R0D8_FOoH;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-k-R#RC80bFRHDbCHRMCW- 
-MRC8DRLFRO	sRNlHDlbCMlC0HN0F#MRHNoMD-#
-CRLoRHM#CCDOs0RNHlRlCbDl0CMNF0HMHR#oDMN#k
VMHO0FoMRCM0_knl_cC58b:0ER0HMCsoC2CRs0MksR0HMCsoCR
H#PHNsNCLDRDPNRH:RMo0CC:sR=;Rj
oLCHRM
RDPNRR:=80CbEc/n;R
RH5VR5b8C0lERFn8Rc>2RR2cURC0EMR
RRNRPD=R:RDPNR4+R;R
RCRM8H
V;RCRs0MksRDPN;M
C8CRo0k_Mlc_n;k
VMHO0FoMRCD0_CFV0P_Csd8.5CEb0RH:RMo0CCRs2skC0sHMRMo0CCHsR#C
Lo
HMRCRs0Mks5b8C0lERFn8Rc
2;CRM8o_C0D0CVFsPC_;d.
MVkOF0HMCRo0C_DVP0FC8s5CEb0RH:RMo0CCRs;lRNG:MRH0CCoss2RCs0kMMRH0CCos#RH
sPNHDNLCNRPDRR:HCM0oRCs:j=R;C
Lo
HMRVRHRC58bR0E-NRlG=R>RRj20MEC
RRRRDPNRR:=80CbERR-l;NG
CRRD
#CRRRRPRND:8=RCEb0;R
RCRM8H
V;RCRs0Mks5DPN2C;
Mo8RCD0_CFV0P;Cs
MVkOF0HMCRo0k_Ml._d5b8C0:ERR0HMCsoC2CRs0MksR0HMCsoCR
H#PHNsNCLDRDPNRH:RMo0CC:sR=;Rj
oLCHRM
RRHV5b8C0<ER=URcR8NMRb8C0>ERR24nRC0EMR
RRPRRN:DR=;R4
CRRMH8RVR;
R0sCkRsMP;ND
8CMR0oC_lMk_;d.
MVkOF0HMCRo0k_Mln_45b8C0:ERR0HMCsoC2CRs0MksR0HMCsoCR
H#PHNsNCLDRDPNRH:RMo0CC:sR=;Rj
oLCHRM
RRHV5b8C0<ER=nR4R8NMRb8C0>ERRRj20MEC
RRRRNRPD=R:R
4;RMRC8VRH;R
RskC0sPMRN
D;CRM8o_C0M_kl4
n;O#FM00NMRlMk_DOCDc_nRH:RMo0CC:sR=CRo0k_Mlc_n5b8C0;E2
MOF#M0N0CRDVP0FCds_.RR:HCM0oRCs:o=RCD0_CFV0P_Csd8.5CEb02O;
F0M#NRM0M_klODCD_Rd.:MRH0CCos=R:R0oC_lMk_5d.D0CVFsPC_2d.;F
OMN#0MD0RCFV0P_Cs4:nRR0HMCsoCRR:=o_C0D0CVFsPC5VDC0CFPs._d,.Rd2O;
F0M#NRM0M_klODCD_R4n:MRH0CCos=R:R0oC_lMk_54nD0CVFsPC_24n;0

$RbCF_k0L_k#0C$b_#ncRRH#NNss$MR5kOl_C_DDn8cRF0IMF,RjR8IH04E-RI8FMR0FjF2RV0R#8F_Do;HO
b0$CkRF0k_L#$_0bdC_.H#R#sRNsRN$5lMk_DOCD._dRI8FMR0FjI,RHE80-84RF0IMF2RjRRFV#_08DHFoO0;
$RbCF_k0L_k#0C$b_#4nRRH#NNss$MR5kOl_C_DD48nRF0IMF,RjR8IH04E-RI8FMR0FjF2RV0R#8F_Do;HO
o#HMRNDs0Fk_#Lk_#ncRF:RkL0_k0#_$_bCn;c#RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-.-R7sRNsRN$F8VRFRk05bHMk00RFsR0H0-#N#0C2H
#oDMNRkIF0k_L#c_n#RR:F_k0L_k#0C$b_#nc;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--.N7Rs$sNRRFV80FkRM5HbRk000FRs#H-0CN0##2
HNoMDFRskL0_kd#_.:#RR0Fk_#Lk_b0$C._d#R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RR.7NNss$VRFRk8F0HR5M0bkRR0F0-sH#00NC
#2#MHoNIDRF_k0L_k#dR.#:kRF0k_L#$_0bdC_.
#;#MHoNsDRF_k0L_k#4Rn#:kRF0k_L#$_0b4C_nR#;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-7R.RsNsNF$RVFR8k50RHkMb0FR0RH0s-N#002C#
o#HMRNDI0Fk_#Lk_#4nRF:RkL0_k0#_$_bC4;n#
o#HMRNDs0Fk__CM#RR:#_08DHFoOC_POs0F5lMk_DOCDc_nRI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-C-RMDNLCV#RF0sRs#H-0CN0#H
#oDMNRkIF0M_C_:#RR8#0_oDFHPO_CFO0sk5MlC_ODnD_cFR8IFM0R;j2
o#HMRNDs0Fk__CMd:.RR8#0_oDFH
O;#MHoNIDRF_k0CdM_.RR:#_08DHFoO#;
HNoMDFRskC0_Mn_4R#:R0D8_FOoH;H
#oDMNRkIF0M_C_R4n:0R#8F_Do;HO
o#HMRNDI_s0C#M_R#:R0D8_FOoH_OPC05FsM_klODCD_Rnc8MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-sRIHR0CCLMNDRC#VRFsCENORIsFRRFV)RqvODCD#H
#oDMNR0Is__CMd:.RR8#0_oDFH
O;#MHoNIDRsC0_Mn_4R#:R0D8_FOoH;H
#oDMNR_HMs_Co#RR:#_08DHFoOC_POs0F58IH04E-RI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RCk#8FR0RosCHC#0sQR7h#R
HNoMDFRsks0_C#o_R#:R0D8_FOoH_OPC05FsI0H8ER-48MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-k-R#RC80sFRC#oH0RCs7amz
o#HMRNDI0Fk_osC_:#RR8#0_oDFHPO_CFO0sH5I8-0E4FR8IFM0R;j2R
RR#MHoNsDRNs8_C#o_R#:R0D8_FOoH_OPC05FsNs88I0H8ER-48MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--k8#CRR0FsHCo#s0CR7q7)H
#oDMNR8IN_osC_:#RR8#0_oDFHPO_CFO0s85N8HsI8-0E4FR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-#RkC08RFCRso0H#CqsR7
7)#MHoNDDRFsI_Ns88_:#RR8#0_oDFHPO_CFO0sR568MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--Ns88R0LH#MRHbRk00)FRqOvRC#DDRR5cL#H0RJsCkCHs8#2
HNoMDFRDIN_I8_8s#RR:#_08DHFoOC_POs0F586RF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-N-R8R8sL#H0RbHMk00RFqR)vCRODRD#5LcRHR0#skCJH8sC2-
-R8CMRD#CCRO0sRNlHDlbCMlC0HN0F#MRHNoMDN#
0H0sLCk0Rs\3NFl_VCV#0:\RRs#0H;Mo
C
Lo
HMRcRzdH:RVsR5Ns88_osC2CRoMNCs0-CR-CRoMNCs0LCRD	FORlsN
RRRRR--QNVR8I8sHE80RO<REOFHCH_I8R0ENH##o'MRj0'RFMRkk8#CR0LH#R
RRjRzRRR:H5VRNs88I0H8ERR=4o2RCsMCN
0CSRRRRIDF_8sN8<sR=jR"jjjjjjjjjjjj"RR&s_N8s5Coj
2;SRRRRIDF_8IN8<sR=jR"jjjjjjjjjjjj"RR&I_N8s5Coj
2;S8CMRMoCC0sNCjRz;R
RR4RzRRR:H5VRNs88I0H8ERR=.o2RCsMCN
0CSFSDIN_s8R8s<"=Rjjjjjjjjjjjj"RR&s_N8s5Co4FR8IFM0R;j2
RSRRFRDIN_I8R8s<"=Rjjjjjjjjjjjj"RR&I_N8s5Co4FR8IFM0R;j2
MSC8CRoMNCs0zCR4R;
RzRR.:RRRRHV58N8s8IH0=ERRRd2oCCMsCN0
DSSFsI_Ns88RR<="jjjjjjjjjjj"RR&s_N8s5Co.FR8IFM0R;j2
RSRRFRDIN_I8R8s<"=Rjjjjjjjjj"jjRI&RNs8_C.o5RI8FMR0Fj
2;S8CMRMoCC0sNC.Rz;R
RRdRzRRR:H5VRNs88I0H8ERR=co2RCsMCN
0CSFSDIN_s8R8s<"=RjjjjjjjjjRj"&NRs8C_soR5d8MFI0jFR2S;
RRRRD_FII8N8s=R<Rj"jjjjjjjjj"RR&I_N8s5CodFR8IFM0R;j2
MSC8CRoMNCs0zCRdR;
RzRRc:RRRRHV58N8s8IH0=ERRR62oCCMsCN0
RSRRFRDIN_s8R8s<"=Rjjjjjjjjj&"RR8sN_osC58cRF0IMF2Rj;R
SRDRRFII_Ns88RR<="jjjjjjjjRj"&NRI8C_soR5c8MFI0jFR2S;
CRM8oCCMsCN0R;zc
RRRRRz6RH:RVNR58I8sHE80Rn=R2CRoMNCs0SC
RRRRD_FIs8N8s=R<Rj"jjjjjjRj"&NRs8C_soR568MFI0jFR2S;
SIDF_8IN8<sR=jR"jjjjj"jjRI&RNs8_C6o5RI8FMR0Fj
2;S8CMRMoCC0sNC6Rz;R
RRnRzRRR:H5VRNs88I0H8ERR=(o2RCsMCN
0CSRRRRIDF_8sN8<sR=jR"jjjjjRj"&NRs8C_soR5n8MFI0jFR2S;
SIDF_8IN8<sR=jR"jjjjjRj"&NRI8C_soR5n8MFI0jFR2S;
CRM8oCCMsCN0R;zn
RRRRRz(RH:RVNR58I8sHE80RU=R2CRoMNCs0SC
RRRRD_FIs8N8s=R<Rj"jjjjj"RR&s_N8s5Co(FR8IFM0R;j2
DSSFII_Ns88RR<="jjjj"jjRI&RNs8_C(o5RI8FMR0Fj
2;S8CMRMoCC0sNC(Rz;R
RRURzRRR:H5VRNs88I0H8ERR=go2RCsMCN
0CSRRRRIDF_8sN8<sR=jR"jjjj"RR&s_N8s5CoUFR8IFM0R;j2
DSSFII_Ns88RR<="jjjjRj"&NRI8C_soR5U8MFI0jFR2S;
CRM8oCCMsCN0R;zU
RRRRRzgRH:RVNR58I8sHE80R4=Rjo2RCsMCN
0CSRRRRIDF_8sN8<sR=jR"j"jjRs&RNs8_Cgo5RI8FMR0Fj
2;SFSDIN_I8R8s<"=Rjjjj"RR&I_N8s5CogFR8IFM0R;j2
MSC8CRoMNCs0zCRgR;
RzRR4RjR:VRHR85N8HsI8R0E=4R42CRoMNCs0SC
RRRRD_FIs8N8s=R<Rj"jj&"RR8sN_osC5R4j8MFI0jFR2S;
SIDF_8IN8<sR=jR"jRj"&NRI8C_soj54RI8FMR0Fj
2;S8CMRMoCC0sNC4RzjR;
RzRR4R4R:VRHR85N8HsI8R0E=.R42CRoMNCs0SC
RRRRD_FIs8N8s=R<Rj"j"RR&s_N8s5Co484RF0IMF2Rj;S
SD_FII8N8s=R<Rj"j"RR&I_N8s5Co484RF0IMF2Rj;C
SMo8RCsMCNR0Cz;44
RRRR.z4RRR:H5VRNs88I0H8ERR=4Rd2oCCMsCN0
RSRRFRDIN_s8R8s<'=Rj&'RR8sN_osC5R4.8MFI0jFR2S;
SIDF_8IN8<sR=jR''RR&I_N8s5Co48.RF0IMF2Rj;C
SMo8RCsMCNR0Cz;4.
RRRRdz4RRR:H5VRNs88I0H8ERR>4Rd2oCCMsCN0
RSRRFRDIN_s8R8s<s=RNs8_C4o5dFR8IFM0R;j2
RSRRFRDIN_I8R8s<I=RNs8_C4o5dFR8IFM0R;j2
MSC8CRoMNCs0zCR4
d;
RRRRR--Q5VR8_HMs2CoRosCHC#0sQR7h#RkHRMoB
piRRRRzR4cRH:RV8R5HsM_CRo2oCCMsCN0
RRRRRRRRFbsO#C#Rp5Bi7,RQRh2LHCoMR
RRRRRRRRRRVRHRp5BiRR='R4'NRM8B'piCMPC002RE
CMRRRRRRRRRRRRRRRRHsM_C<oR="R5jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"RR&72Qh;R
RRRRRRRRRRMRC8VRH;R
RRRRRRMRC8sRbF#OC#S;
CRM8oCCMsCN0Rcz4;R
RR4Rz6:RRRRHV50MFRM8H_osC2CRoMNCs0RC
RRRRRRRRRHRRMC_so=R<Rj5"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jjR7&RQ;h2
MSC8CRoMNCs0zCR4
6;
RRRRR--Q5VRsk8F0C_sos2RC#oH0RCs)m_7zkaR#oHMRm)_B
piRRRRzs4n80FkRRR:H5VRsk8F0C_soo2RCsMCN
0CRRRRRRRRbOsFCR##5m)_B,piRksF0C_soL2RCMoH
RRRRRRRRRRRRRHV5m)_BRpi=4R''MRN8_R)miBp'CCPMR020MEC
RRRRRRRRRRRRRRRR7)_mRza<s=RF_k0s4Co;R
RRRRRRRRRRMRC8VRH;R
RRRRRRMRC8sRbF#OC#R;
RRRRRCRRMo8RCsMCNR0Czs4n80Fk;R
RR4Rz(Fs8kR0R:VRHRF5M08RsF_k0s2CoRMoCC0sNCR
RRRRRRRRRR_R)7amzRR<=s0Fk_osC4S;
CRM8oCCMsCN0R(z4sk8F0
;
Snz4Ik8F0:RRRRHV5FI8ks0_CRo2oCCMsCN0
RRRRRRRRFbsO#C#R_5WmiBp,FRIks0_CRo2LHCoMR
RRRRRRRRRRVRHR_5WmiBpR'=R4N'RMW8R_pmBiP'CC2M0RC0EMR
RRRRRRRRRRRRRR_RW7amzRR<=I0Fk_osC58IH04E-RI8FMR0Fj
2;RRRRRRRRRRRRCRM8H
V;RRRRRRRRCRM8bOsFC;##
RRRRRRRR8CMRMoCC0sNC4RznFI8k
0;RRRRzI4(80FkRRR:H5VRMRF0Ik8F0C_soo2RCsMCN
0CRRRRRRRRRRRRWm_7z<aR=FRIks0_CIo5HE80-84RF0IMF2Rj;C
SMo8RCsMCNR0CzI4(80Fk;R

R-RR-VRQRN5s8_8ss2CoRosCHC#0sqR)7R7)kM#HoBRmpRi
RzRR4RnsRH:RVsR5Ns88_osC2CRoMNCs0-C
-RRRRRRRRFbsO#C#RB5mpRi,)7q7)L2RCMoH
R--RRRRRRRRRHRRVmR5BRpi=4R''MRN8BRmpCi'P0CM2ER0C-M
-RRRRRRRRRRRRRRRR8sN_osCRR<=)7q7)85N8HsI8-0E4FR8IFM0R;j2
R--RRRRRRRRRCRRMH8RV-;
-RRRRRRRR8CMRFbsO#C#;-
-S8CMRMoCC0sNC4Rzn
s;-R-RR4Rz(:sRRRHV50MFR8sN8ss_CRo2oCCMsCN0
RRRRRRRRRRRR8sN_osCRR<=)7q7)S;
CRM8oCCMsCN0Rnz4s
;
SR--Q5VRI8N8sC_sos2RC#oH0RCsW7q7)#RkHRMoWB_mpRi
RzRR4RnIRH:RVIR5Ns88_osC2CRoMNCs0RC
RRRRRbRRsCFO#5#RB,piR7Wq7R)2LHCoMR
RRRRRRRRRRVRHRp5BiRR='R4'NRM8B'piCMPC002RE
CMRRRRRRRRRRRRRRRRI_N8sRCo<W=Rq)7758N8s8IH04E-RI8FMR0Fj
2;RRRRRRRRRRRRCRM8H
V;RRRRRRRRCRM8bOsFC;##
MSC8CRoMNCs0zCR4;nI
RRRR(z4IRR:H5VRMRF0I8N8sC_soo2RCsMCN
0CRRRRRRRRRRRRI_N8sRCo<W=Rq)77;C
SMo8RCsMCNR0CzI4(;R

R-RR-GR 0RsNDHFoOFRVskR7NbDRFRs0OCN#
sSzC:oRRFbsO#C#5iBp2CRLo
HMSHRRVBR5p i'ea hR8NMRiBpR'=R4R'20MEC
RSRRh7Q_b0lRR<=7;Qh
RSRR7)q70)_l<bR=qR)7;7)
RSRR7Wq70)_l<bR=qRW7;7)
RSRR_W 0Rlb<W=R S;
RMRC8VRH;C
SMb8RsCFO#
#;
-S-RRQV)8CNR8q8s#C#RW=RsCH0R8q8s#C#,$RLb#N#Rh7QRR0FFbk0kH0RV RWRRH#CLMND
C8SkzlGRR:bOsFC5##W0 _lRb,)7q7)l_0bW,Rq)77_b0l,QR7hl_0bs,RF_k0s2Co
RSRLHCoMR
SRHRRVWR5q)77_b0lR)=Rq)77_b0lR8NMR_W 0Rlb=4R''02RE
CMSRSRs0Fk_osC4=R<Rh7Q_b0l;S
SCCD#
RSSRksF0C_so<4R=FRsks0_CIo5HE80-84RF0IMF2Rj;S
SCRM8H
V;S8CMRFbsO#C#;R
SR
RRRRRR-t-RCsMCNR0C0REC)RqvODCD#MRN8CR#D0CORoDFHVORF)sRq4vAn4_1_
14SUz4RH:RVOR5EOFHCH_I8R0E=2R4RMoCC0sNCR
RRzRS4:gRRsVFRHHRM8R5CEb0_lMk_DOCD-#RRR428MFI0jFRRMoCC0sNC-
S-VRQR85N8HsI8R0E>cR42CRMC08RFsROCCN0RHIs0CCRMDNLCMRN8kRF00bkRNCMLRDC#CCDOD0RFOoH
RRRRRRRR.SzjRR:H5VRNs88I0H8ERR>4Rc2oCCMsCN0
-S-RGVHRsVFRDONDdR4U,U(RD#CCRO0F0VRs0H#NR0CMRF0LMCHoCRso0H#C8sC
SSSSksF0M_C5RH2<'=R4I'RERCM57)q70)_lNb58I8sHE80-84RF0IMFcR42RR=HC2RDR#C';j'
SSSSkIF0M_C5RH2<'=R4I'RERCM58IN_osC58N8s8IH04E-RI8FMR0F4Rc2=2RHR#CDCjR''R;
RRRRRRRRRRRRRIRRsC0_M25HRR<=WI RERCM58IN_osC58N8s8IH04E-RI8FMR0F4Rc2=2RHR#CDCjR''R;
RRRRRSRRCRM8oCCMsCN0Rjz.;-
S-VRQR85N8HsI8R0E<4=RcM2RFsRIHR0CCLMNDFCRskRF00bkRNCMLRDC#CCDOD0RFOoHRCMC8
C8RRSRRzRS.:4RRRHV58N8s8IH0<ER=cR42CRoMNCs0SC
SsSSF_k0CHM52=R<R''4;S
SSFSIkC0_M25HRR<=';4'
RRRRRRRRRRRRRRRR0Is_5CMH<2R= RW;R
RRRRRRCRSMo8RCsMCNR0Cz;.4
-S-RMtCC0sNCER0CqR)vCRODRD#NRM80-sH#00NCR#
RRRRRSRRzR..:FRVsRR[H5MRI0H8Ek_MlC_ODRD#-2R4RI8FMR0FjCRoMNCs0RC
RRRRRRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)RAq4v_ncdUXR47:NRDLRCDH"#RW
";RRRRRRRRRRRRRRRRLHCoMR
RRRRRRRRRRARS)_qv4Undc7X4R):Rq4vAn4_1_
14SRRRRRRRRRRRRsbF0NRlb7R5Qjq52>R=R_HMs5Co[R2,q)77q>R=RIDF_8IN84s5dFR8IFM0R,j2RA7QRR=>",j"R7q7)=AR>FRDIN_s858s48dRF0IMF2Rj,S
SShS q>R=R''4,1R1)=qR>jR''W,R =qR>sRI0M_C5,H2RiBpq>R=RiBp,hR A>R=R''4,1R1)=AR>jR''W,R =AR>jR''B,RpRiA=B>Rp
i,SRSSR7RRmjq52>R=RkIF0k_L#H45,,[2RA7m5Rj2=s>RF_k0L4k#5[H,2
2;
RRRRRRRRRRRRRRRRksF0C_so25[RR<=s0Fk_#Lk4,5H[I2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
SSSSkIF0C_so25[RR<=I0Fk_#Lk4,5HKI2RERCM5kIF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRMSC8CRoMNCs0zCR.
.;RRRRRMSC8CRoMNCs0zCR4
g;RRRRCRM8oCCMsCN0RUz4;RRRRR
RRRRR
RRRRR--tCCMsCN0RC0ERv)qRDOCDN#RM#8RCODC0FRDoRHOVRFs)Aqv41n_.._1
.SzdRR:H5VROHEFOIC_HE80R.=R2CRoMNCs0RC
RSRRzR.c:FRVsRRHH5MR80CbEk_MlC_ODRD#-2R4RI8FMR0FjCRoMNCs0SC
-Q-RVNR58I8sHE80R4>RdM2RCRC80OFRs0CNCsRIHR0CCLMNDNCRMF8Rkk0b0MRCNCLDRD#CCRO0DHFoOR
RRRRRRzRS.:6RRRHV58N8s8IH0>ERR24dRMoCC0sNC-
S-HRVGFRVsNROD4DRd(UU,CR#D0CORRFV0#sH0CN0R0MFRHLCMsoRC#oH0CCs8R
RRRRRRRRRRRRRRFRskC0_M25HRR<='R4'IMECRq5)7_7)05lbNs88I0H8ER-48MFI04FRd=2RRRH2CCD#R''j;S
SSFSIkC0_M25HRR<='R4'IMECRN5I8C_so85N8HsI8-0E4FR8IFM0R24dRH=R2DRC#'CRj
';RRRRRRRRRRRRRRRRI_s0CHM52=R<RRW IMECRN5I8C_so85N8HsI8-0E4FR8IFM0R24dRH=R2DRC#'CRj
';RRRRRRRRS8CMRMoCC0sNC.Rz6S;
-Q-RVNR58I8sHE80RR<=4Rd2MIFRsCH0RNCMLRDCFFsRkk0b0MRCNCLDRD#CCRO0DHFoOCRMC88C
RRSRSRRzR.n:VRHR85N8HsI8R0E<4=Rdo2RCsMCN
0CSRRRRRRRRRRRRksF0M_C5RH2<'=R4
';SSSSI0Fk_5CMH<2R=4R''R;
RRRRRRRRRRRRRIRRsC0_M25HRR<=W
 ;RRRRRRRRS8CMRMoCC0sNC.RznS;
-t-RCsMCNR0C0REC)RqvODCD#MRN8sR0H0-#N#0C
RRRRRRRR.Sz(RR:VRFs[MRHRH5I8_0EM_klODCD#RR-482RF0IMFRRjoCCMsCN0
RRRRRRRRRRRRRRRR0N0skHL0\CR3lsN_VFV#\C0RRFVAv)q_gU4.7X.RD:RNDLCRRH#";W"
RRRRRRRRRRRRRRRRoLCHRM
RRRRRRRRRSRRAv)q_gU4.7X.R):Rq4vAn._1_
1.SRRRRRRRRRRRRsbF0NRlb7R5Q=qR>MRH_osC5[.*+84RF0IMF*R.[R2,q)77q>R=RIDF_8IN84s5.FR8IFM0R,j2RA7QRR=>""jj,7Rq7R)A=D>RFsI_Ns885R4.8MFI0jFR2S,
SRSRRhR q>R=R''4,1R1)=qR>jR''W,R =qR>sRI0M_C5,H2RiBpq>R=RiBp,hR A>R=R''4,1R1)=AR>jR''W,R =AR>jR''B,RpRiA=B>Rp
i,SRSSR7RRm4q52>R=RkIF0k_L#H.5,[.*+,42Rq7m5Rj2=I>RF_k0L.k#5.H,*,[2RA7m5R42=s>RF_k0L.k#5.H,*4[+27,RmjA52>R=RksF0k_L#H.5,*R.[;22
RRRRRRRRRRRRRRRRksF0C_so*5.[<2R=FRskL0_k5#.H*,.[I2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRksF0C_so*5.[2+4RR<=s0Fk_#Lk.,5H.+*[4I2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
SSSSkIF0C_so*5.[<2R=FRIkL0_k5#.H*,.[I2RERCM5kIF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRkIF0C_so*5.[2+4RR<=I0Fk_#Lk.,5H.+*[4I2RERCM5kIF0M_C5RH2=4R''C2RDR#C';Z'
R
RRRRRRCRSMo8RCsMCNR0Cz;.(
RRRRCRSMo8RCsMCNR0Cz;.c
RRRR8CMRMoCC0sNC.RzdR;R
R
SR-RR-CRtMNCs00CRE)CRqOvRC#DDR8NMRD#CCRO0DHFoOFRVsqR)vnA4__1c1Sc
zR.U:VRHRE5OFCHO_8IH0=ERRRc2oCCMsCN0
RRRR.SzgRR:VRFsHMRHRC58b_0EM_klODCD#RR-482RF0IMFRRjoCCMsCN0
-S-RRQV58N8s8IH0>ERR24.RCMC8FR0RCOsNR0CI0sHCMRCNCLDR8NMR0FkbRk0CLMND#CRCODC0FRDo
HORRRRRRRRSjzdRH:RVNR58I8sHE80R4>R.o2RCsMCN
0CSR--VRHGVRFsODNDRU4dUR(,#CCDOF0RVsR0HN#00MCRFL0RCoHMRosCHC#0s
C8RRRRRRRRRRRRRRRRs0Fk_5CMH<2R=4R''ERIC5MR)7q7)l_0b85N8HsI8-0E4FR8IFM0R24.RH=R2DRC#'CRj
';SSSSI0Fk_5CMH<2R=4R''ERIC5MRI_N8s5CoNs88I0H8ER-48MFI04FR.-2RRRH2CCD#R''j;R
RRRRRRRRRRRRRRsRI0M_C5RH2<W=R ERIC5MRI_N8s5CoNs88I0H8ER-48MFI04FR.=2RRRH2CCD#R''j;R
RRRRRRCRSMo8RCsMCNR0Cz;dj
-S-RRQV58N8s8IH0<ER=.R42FRMRHIs0CCRMDNLCsRFR0FkbRk0CLMND#CRCODC0FRDoRHOM8CCCR8
SRRRRdSz4RR:H5VRNs88I0H8E=R<R24.RMoCC0sNCS
SSFSskC0_M25HRR<=';4'
SSSSkIF0M_C5RH2<'=R4
';RRRRRRRRRRRRRRRRI_s0CHM52=R<R;W 
RRRRRRRRMSC8CRoMNCs0zCRd
4;SR--tCCMsCN0RC0ERv)qRDOCDN#RM08Rs#H-0CN0#R
RRRRRRzRSd:.RRsVFRH[RMIR5HE80_lMk_DOCD-#RRR428MFI0jFRRMoCC0sNCR
RRRRRRRRRRRRRR0RN0LsHkR0C\N3slV_FV0#C\VRFRqA)vj_cgcnX7RR:DCNLD#RHR""W;R
RRRRRRRRRRRRRRCRLo
HMRRRRRRRRRRRRSqA)vj_cgcnX7RR:)Aqv41n_cc_1
RSRRRRRRRRRRFRbsl0RN5bR7RQq=H>RMC_so*5c[R+d8MFI0cFR*,[2R7q7)=qR>FRDIN_I858s484RF0IMF2Rj,QR7A>R=Rj"jj,j"R7q7)=AR>FRDIN_s858s484RF0IMF2Rj,S
SShS q>R=R''4,1R1)=qR>jR''W,R =qR>sRI0M_C5,H2RiBpq>R=RiBp,hR A>R=R''4,1R1)=AR>jR''W,R =AR>jR''B,RpRiA=B>Rp
i,SSSS75mqd=2R>FRIkL0_k5#cHc,R*d[+2
,RSSSS75mq.=2R>FRIkL0_k5#cH*,c[2+.,SR
S7SSm4q52>R=RkIF0k_L#Hc5,[c*+,42RS
SSmS7q25jRR=>I0Fk_#Lkc,5HR[c*2S,
S7SSmdA52>R=RksF0k_L#Hc5,*Rc[2+d,SR
S7SSm.A52>R=RksF0k_L#Hc5,[c*+,.2RS
SSmS7A254RR=>s0Fk_#Lkc,5Hc+*[4R2,
SSSSA7m5Rj2=s>RF_k0Lck#5RH,c2*[2S;
SsSSF_k0s5Coc2*[RR<=s0Fk_#Lkc,5Hc2*[RCIEMsR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRsRRF_k0s5Coc+*[4<2R=FRskL0_k5#cH*,c[2+4RCIEMsR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRsRRF_k0s5Coc+*[.<2R=FRskL0_k5#cH*,c[2+.RCIEMsR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRsRRF_k0s5Coc+*[d<2R=FRskL0_k5#cH*,c[2+dRCIEMsR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRIRRF_k0s5Coc2*[RR<=I0Fk_#Lkc,5Hc2*[RCIEMIR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRIRRF_k0s5Coc+*[4<2R=FRIkL0_k5#cH*,c[2+4RCIEMIR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRIRRF_k0s5Coc+*[.<2R=FRIkL0_k5#cH*,c[2+.RCIEMIR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRIRRF_k0s5Coc+*[d<2R=FRIkL0_k5#cH*,c[2+dRCIEMIR5F_k0CHM52RR='24'R#CDCZR''
;
RRRRRRRRS8CMRMoCC0sNCdRz.R;
RRRRS8CMRMoCC0sNC.RzgR;
RCRRMo8RCsMCNR0Cz;.U
R
SR-RR-CRtMNCs00CRE)CRqOvRC#DDR8NMRD#CCRO0DHFoOFRVsqR)vnA4__1g1Sg
zRdd:VRHRE5OFCHO_8IH0=ERRRg2oCCMsCN0
RRRRdSzcRR:VRFsHMRHRC58b_0EM_klODCD#RR-482RF0IMFRRjoCCMsCN0
-S-RRQV58N8s8IH0>ERR244RCMC8FR0RCOsNR0CI0sHCMRCNCLDR8NMR0FkbRk0CLMND#CRCODC0FRDo
HORRRRRRRRS6zdRH:RVNR58I8sHE80R4>R4o2RCsMCN
0CSR--VRHGVRFsODNDRU4dUR(,#CCDOF0RVsR0HN#00MCRFL0RCoHMRosCHC#0s
C8RRRRRRRRRRRRRRRRs0Fk_5CMH<2R=4R''ERIC5MR)7q7)l_0b85N8HsI8-0E4FR8IFM0R244RH=R2DRC#'CRj
';SSSSI0Fk_5CMH<2R=4R''ERIC5MRI_N8s5CoNs88I0H8ER-48MFI04FR4=2RRRH2CCD#R''j;R
RRRRRRRRRRRRRRsRI0M_C5RH2<W=R ERIC5MRI_N8s5CoNs88I0H8ER-48MFI04FR4=2RRRH2CCD#R''j;R
RRRRRRCRSMo8RCsMCNR0Cz;d6
-S-RRQV58N8s8IH0<ER=4R42FRMRHIs0CCRMDNLCsRFR0FkbRk0CLMND#CRCODC0FRDoRHOM8CCCR8
SRRRRdSznRR:H5VRNs88I0H8E=R<R244RMoCC0sNCR
SRRRRRRRRRsRRF_k0CHM52=R<R''4;S
SSFSIkC0_M25HRR<=';4'
RRRRRRRRRRRRRRRR0Is_5CMH<2R= RW;R
RRRRRRCRSMo8RCsMCNR0Cz;dn
-S-RMtCC0sNCER0CqR)vCRODRD#NRM80-sH#00NCR#
RRRRRSRRzRd(:FRVsRR[H5MRI0H8Ek_MlC_ODRD#-2R4RI8FMR0FjCRoMNCs0RC
RRRRRRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)RAq.v_jXcUU:7RRLDNCHDR#WR""R;
RRRRRRRRRRRRRLRRCMoH
RRRRRRRRRRRR)SAq.v_jXcUU:7RRv)qA_4n11g_gR
RRRRRRRRRRRRRRRRRb0FsRblNRQ57q>R=R_HMs5Cog+*[(FR8IFM0R[g*2q,R7q7)RR=>D_FII8N8sj54RI8FMR0FjR2,7RQA=">Rjjjjjjjj"q,R7A7)RR=>D_FIs8N8sj54RI8FMR0Fj
2,RRRRRRRRRRRRRRRRRRRRRRRRRRRR Rhq='>R4R',1q1)RR=>',j'RqW RR=>I_s0CHM52B,RpRiq=B>RpRi, RhA='>R4R',1A1)RR=>',j'RAW RR=>',j'RiBpA>R=RiBp,RR
RRRRRRRRRRRRRRRRRRRRRRRRR7RRm(q52>R=RkIF0k_L#HU5,[U*+,(2RR
RRRRRRRRRRRRRRRRRRRRRRRRRRmR7q25nRR=>I0Fk_#LkU,5HU+*[nR2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRq7m5R62=I>RF_k0LUk#5UH,*6[+2
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mqc=2R>FRIkL0_k5#UH*,U[2+c,RR
RRRRRRRRRRRRRRRRRRRRRRRRR7RRmdq52>R=RkIF0k_L#HU5,[U*+,d2RR
RRRRRRRRRRRRRRRRRRRRRRRRRRmR7q25.RR=>I0Fk_#LkU,5HU+*[.R2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRq7m5R42=I>RF_k0LUk#5UH,*4[+2
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mqj=2R>FRIkL0_k5#UH*,U[R2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRA7m5R(2=s>RF_k0LUk#5UH,*([+2
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mAn=2R>FRskL0_k5#UH*,U[2+n,RR
RRRRRRRRRRRRRRRRRRRRRRRRR7RRm6A52>R=RksF0k_L#HU5,[U*+,62RR
RRRRRRRRRRRRRRRRRRRRRRRRRRmR7A25cRR=>s0Fk_#LkU,5HU+*[cR2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRA7m5Rd2=s>RF_k0LUk#5UH,*d[+2
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mA.=2R>FRskL0_k5#UH*,U[2+.,RR
RRRRRRRRRRRRRRRRRRRRRRRRR7RRm4A52>R=RksF0k_L#HU5,[U*+,42RR
RRRRRRRRRRRRRRRRRRRRRRRRRRmR7A25jRR=>s0Fk_#LkU,5HU2*[,RR
RRRRRRRRRRRRRRRRRRRRRRRRR7RRQ5uqj=2R>MRH_osC5[g*+,U2Ru7QA>R=R""j,R
RRRRRRRRRRRRRRRRRRRRRRRRRRmR7ujq52>R=RNIbs$H0_#LkU,5H[R2,7Amu5Rj2=s>RbHNs0L$_k5#UH2,[2R;
RRRRRRRRRRRRRsRRF_k0s5Cog2*[RR<=s0Fk_#LkU,5HU2*[RCIEMsR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRsRRF_k0s5Cog+*[4<2R=FRskL0_k5#UH*,U[2+4RCIEMsR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRsRRF_k0s5Cog+*[.<2R=FRskL0_k5#UH*,U[2+.RCIEMsR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRsRRF_k0s5Cog+*[d<2R=FRskL0_k5#UH*,U[2+dRCIEMsR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRsRRF_k0s5Cog+*[c<2R=FRskL0_k5#UH*,U[2+cRCIEMsR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRsRRF_k0s5Cog+*[6<2R=FRskL0_k5#UH*,U[2+6RCIEMsR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRsRRF_k0s5Cog+*[n<2R=FRskL0_k5#UH*,U[2+nRCIEMsR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRsRRF_k0s5Cog+*[(<2R=FRskL0_k5#UH*,U[2+(RCIEMsR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRsRRF_k0s5Cog+*[U<2R=bRsN0sH$k_L#HU5,R[2IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRFRIks0_Cgo5*R[2<I=RF_k0LUk#5UH,*R[2IMECRF5IkC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRFRIks0_Cgo5*4[+2=R<RkIF0k_L#HU5,[U*+R42IMECRF5IkC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRFRIks0_Cgo5*.[+2=R<RkIF0k_L#HU5,[U*+R.2IMECRF5IkC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRFRIks0_Cgo5*d[+2=R<RkIF0k_L#HU5,[U*+Rd2IMECRF5IkC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRFRIks0_Cgo5*c[+2=R<RkIF0k_L#HU5,[U*+Rc2IMECRF5IkC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRFRIks0_Cgo5*6[+2=R<RkIF0k_L#HU5,[U*+R62IMECRF5IkC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRFRIks0_Cgo5*n[+2=R<RkIF0k_L#HU5,[U*+Rn2IMECRF5IkC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRFRIks0_Cgo5*([+2=R<RkIF0k_L#HU5,[U*+R(2IMECRF5IkC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRFRIks0_Cgo5*U[+2=R<RNIbs$H0_#LkU,5H[I2RERCM5kIF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRMSC8CRoMNCs0zCRd
(;RRRRRMSC8CRoMNCs0zCRd
c;RRRRCRM8oCCMsCN0Rdzd;S

RRRR-t-RCsMCNR0C0REC)RqvODCD#MRN8CR#D0CORoDFHVORF)sRq4vAn4_1U4_1Uz
Sd:URRRHV5FOEH_OCI0H8ERR=4RU2oCCMsCN0
RRRRdSzgRR:VRFsHMRHRC58b_0EM_klODCD#RR-482RF0IMFRRjoCCMsCN0
-S-RRQV58N8s8IH0>ERR24jRCMC8FR0RCOsNR0CI0sHCMRCNCLDR8NMR0FkbRk0CLMND#CRCODC0FRDo
HORRRRRRRRSjzcRH:RVNR58I8sHE80R4>Rjo2RCsMCN
0CSR--VRHGVRFsODNDRU4dUR(,#CCDOF0RVsR0HN#00MCRFL0RCoHMRosCHC#0s
C8RRRRRRRRRRRRRRRRs0Fk_5CMH<2R=4R''ERIC5MR)7q7)l_0b85N8HsI8-0E4FR8IFM0R24jRH=R2DRC#'CRj
';SSSSI0Fk_5CMH<2R=4R''ERIC5MRI_N8s5CoNs88I0H8ER-48MFI04FRj=2RR2HRR#CDCjR''R;
RRRRRRRRRRRRRIRRsC0_M25HRR<=WI RERCM58IN_osC58N8s8IH04E-RI8FMR0F4Rj2=2RHR#CDCjR''R;
RRRRRSRRCRM8oCCMsCN0Rjzc;-
S-VRQR85N8HsI8R0E<4=RjM2RFsRIHR0CCLMNDFCRskRF00bkRNCMLRDC#CCDOD0RFOoHRCMC8
C8RRSRRzRSc:4RRRHV58N8s8IH0<ER=jR42CRoMNCs0SC
RRRRRRRRRRRRs0Fk_5CMH<2R=4R''S;
SISSF_k0CHM52=R<R''4;R
RRRRRRRRRRRRRRsRI0M_C5RH2<W=R R;
RRRRRSRRCRM8oCCMsCN0R4zc;-
S-CRtMNCs00CRE)CRqOvRC#DDR8NMRH0s-N#00
C#RRRRRRRRS.zcRV:RF[sRRRHM58IH0ME_kOl_C#DDR4-R2FR8IFM0RojRCsMCN
0CRRRRRRRRRRRRRRRRNs00H0LkC3R\s_NlF#VVCR0\FAVR)_qv4cj.X74nRD:RNDLCRRH#";W"
RRRRRRRRRRRRRRRRoLCHRM
RRRRRRRRRSRRAv)q_.4jcnX47RR:)Aqv41n_41U_4RU
RRRRRRRRRRRRRRRRRsbF0NRlb7R5Q=qR>MRH_osC5*4U[6+4RI8FMR0F4[U*2q,R7q7)RR=>D_FII8N8sR5g8MFI0jFR27,RQ=AR>jR"jjjjjjjjjjjjj"jj,7Rq7R)A=D>RFsI_Ns8858gRF0IMF2Rj,R
RRRRRRRRRRRRRRRRRRRRRRRRRRhR q>R=R''4,1R1)=qR>jR''W,R =qR>sRI0M_C5,H2RiBpq>R=RiBp,hR A>R=R''4,1R1)=AR>jR''W,R =AR>jR''B,RpRiA=B>RpRi,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRq7m5246RR=>I0Fk_#Lk4Hn5,*4n[6+42
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mq4Rc2=I>RF_k0L4k#n,5H4[n*+24c,RR
RRRRRRRRRRRRRRRRRRRRRRRRR7RRm4q5d=2R>FRIkL0_kn#454H,n+*[4,d2RR
RRRRRRRRRRRRRRRRRRRRRRRRRRmR7q.542>R=RkIF0k_L#54nHn,4*4[+.R2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRq7m5244RR=>I0Fk_#Lk4Hn5,*4n[4+42
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mq4Rj2=I>RF_k0L4k#n,5H4[n*+24j,RR
RRRRRRRRRRRRRRRRRRRRRRRRR7RRmgq52>R=RkIF0k_L#54nHn,4*g[+2
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mqU=2R>FRIkL0_kn#454H,n+*[UR2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRq7m5R(2=I>RF_k0L4k#n,5H4[n*+,(2RR
RRRRRRRRRRRRRRRRRRRRRRRRRRmR7q25nRR=>I0Fk_#Lk4Hn5,*4n[2+n,RR
RRRRRRRRRRRRRRRRRRRRRRRRR7RRm6q52>R=RkIF0k_L#54nHn,4*6[+2
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mqc=2R>FRIkL0_kn#454H,n+*[cR2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRq7m5Rd2=I>RF_k0L4k#n,5H4[n*+,d2RR
RRRRRRRRRRRRRRRRRRRRRRRRRRmR7q25.RR=>I0Fk_#Lk4Hn5,*4n[2+.,RR
RRRRRRRRRRRRRRRRRRRRRRRRR7RRm4q52>R=RkIF0k_L#54nHn,4*4[+2
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mqj=2R>FRIkL0_kn#454H,n2*[,RR
RRRRRRRRRRRRRRRRRRRRRRRRR7RRm4A56=2R>FRskL0_kn#454H,n+*[4,62RR
RRRRRRRRRRRRRRRRRRRRRRRRRRmR7Ac542>R=RksF0k_L#54nHn,4*4[+cR2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRA7m524dRR=>s0Fk_#Lk4Hn5,*4n[d+42
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mA4R.2=s>RF_k0L4k#n,5H4[n*+24.,RR
RRRRRRRRRRRRRRRRRRRRRRRRR7RRm4A54=2R>FRskL0_kn#454H,n+*[4,42RR
RRRRRRRRRRRRRRRRRRRRRRRRRRmR7Aj542>R=RksF0k_L#54nHn,4*4[+jR2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRA7m5Rg2=s>RF_k0L4k#n,5H4[n*+,g2RR
RRRRRRRRRRRRRRRRRRRRRRRRRRmR7A25URR=>s0Fk_#Lk4Hn5,*4n[2+U,RR
RRRRRRRRRRRRRRRRRRRRRRRRR7RRm(A52>R=RksF0k_L#54nHn,4*([+2
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mAn=2R>FRskL0_kn#454H,n+*[nR2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRA7m5R62=s>RF_k0L4k#n,5H4[n*+,62RR
RRRRRRRRRRRRRRRRRRRRRRRRRRmR7A25cRR=>s0Fk_#Lk4Hn5,*4n[2+c,RR
RRRRRRRRRRRRRRRRRRRRRRRRR7RRmdA52>R=RksF0k_L#54nHn,4*d[+2
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mA.=2R>FRskL0_kn#454H,n+*[.R2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRA7m5R42=s>RF_k0L4k#n,5H4[n*+,42RR
RRRRRRRRRRRRRRRRRRRRRRRRRRmR7A25jRR=>s0Fk_#Lk4Hn5,*4n[R2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRu7Qq>R=R_HMs5Co4[U*+R4(8MFI04FRU+*[4,n2Ru7QA>R=Rj"j"R,
RRRRRRRRRRRRRRRRRRRRRRRRR7RRm5uq4=2R>bRIN0sH$k_L#54nH*,.[2+4,mR7ujq52>R=RNIbs$H0_#Lk4Hn5,[.*2R,
RRRRRRRRRRRRRRRRRRRRRRRRR7RRm5uA4=2R>bRsN0sH$k_L#54nH*,.[2+4,mR7ujA52>R=RNsbs$H0_#Lk4Hn5,[.*2
2;RRRRRRRRRRRRRRRRs0Fk_osC5*4U[<2R=FRskL0_kn#454H,n2*[RCIEMsR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRsRRF_k0s5Co4[U*+R42<s=RF_k0L4k#n,5H4[n*+R42IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRFRsks0_C4o5U+*[.<2R=FRskL0_kn#454H,n+*[.I2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRksF0C_soU54*d[+2=R<RksF0k_L#54nHn,4*d[+2ERIC5MRs0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRs0Fk_osC5*4U[2+cRR<=s0Fk_#Lk4Hn5,*4n[2+cRCIEMsR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRsRRF_k0s5Co4[U*+R62<s=RF_k0L4k#n,5H4[n*+R62IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRFRsks0_C4o5U+*[n<2R=FRskL0_kn#454H,n+*[nI2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRksF0C_soU54*([+2=R<RksF0k_L#54nHn,4*([+2ERIC5MRs0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRs0Fk_osC5*4U[2+URR<=s0Fk_#Lk4Hn5,*4n[2+URCIEMsR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRsRRF_k0s5Co4[U*+Rg2<s=RF_k0L4k#n,5H4[n*+Rg2IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRFRsks0_C4o5U+*[4Rj2<s=RF_k0L4k#n,5H4[n*+24jRCIEMsR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRsRRF_k0s5Co4[U*+244RR<=s0Fk_#Lk4Hn5,*4n[4+42ERIC5MRs0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRs0Fk_osC5*4U[.+42=R<RksF0k_L#54nHn,4*4[+.I2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRksF0C_soU54*4[+d<2R=FRskL0_kn#454H,n+*[4Rd2IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRFRsks0_C4o5U+*[4Rc2<s=RF_k0L4k#n,5H4[n*+24cRCIEMsR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRsRRF_k0s5Co4[U*+246RR<=s0Fk_#Lk4Hn5,*4n[6+42ERIC5MRs0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRs0Fk_osC5*4U[n+42=R<RNsbs$H0_#Lk4Hn5,[.*2ERIC5MRs0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRs0Fk_osC5*4U[(+42=R<RNsbs$H0_#Lk4Hn5,[.*+R42IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R

RRRRRRRRRRRRRIRRF_k0s5Co4[U*2=R<RkIF0k_L#54nHn,4*R[2IMECRF5IkC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRFRIks0_C4o5U+*[4<2R=FRIkL0_kn#454H,n+*[4I2RERCM5kIF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRkIF0C_soU54*.[+2=R<RkIF0k_L#54nHn,4*.[+2ERIC5MRI0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRI0Fk_osC5*4U[2+dRR<=I0Fk_#Lk4Hn5,*4n[2+dRCIEMIR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRIRRF_k0s5Co4[U*+Rc2<I=RF_k0L4k#n,5H4[n*+Rc2IMECRF5IkC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRFRIks0_C4o5U+*[6<2R=FRIkL0_kn#454H,n+*[6I2RERCM5kIF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRkIF0C_soU54*n[+2=R<RkIF0k_L#54nHn,4*n[+2ERIC5MRI0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRI0Fk_osC5*4U[2+(RR<=I0Fk_#Lk4Hn5,*4n[2+(RCIEMIR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRIRRF_k0s5Co4[U*+RU2<I=RF_k0L4k#n,5H4[n*+RU2IMECRF5IkC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRFRIks0_C4o5U+*[g<2R=FRIkL0_kn#454H,n+*[gI2RERCM5kIF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRkIF0C_soU54*4[+j<2R=FRIkL0_kn#454H,n+*[4Rj2IMECRF5IkC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRFRIks0_C4o5U+*[4R42<I=RF_k0L4k#n,5H4[n*+244RCIEMIR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRIRRF_k0s5Co4[U*+24.RR<=I0Fk_#Lk4Hn5,*4n[.+42ERIC5MRI0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRI0Fk_osC5*4U[d+42=R<RkIF0k_L#54nHn,4*4[+dI2RERCM5kIF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRkIF0C_soU54*4[+c<2R=FRIkL0_kn#454H,n+*[4Rc2IMECRF5IkC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRFRIks0_C4o5U+*[4R62<I=RF_k0L4k#n,5H4[n*+246RCIEMIR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRIRRF_k0s5Co4[U*+24nRR<=IsbNH_0$L4k#n,5H.2*[RCIEMIR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRIRRF_k0s5Co4[U*+24(RR<=IsbNH_0$L4k#n,5H.+*[4I2RERCM5kIF0M_C5RH2=4R''C2RDR#C';Z'
R
RRRRRRCRSMo8RCsMCNR0Cz;c.
RRRRCRSMo8RCsMCNR0Cz;dg
RRRR8CMRMoCC0sNCdRzU
;
SRRRRR--tCCMsCN0RC0ERv)qRDOCDN#RM#8RCODC0FRDoRHOVRFs)Aqv41n_d1n_dSn
zNdURH:RVOR5EOFHCH_I8R0E=nRd2CRoMNCs0SC
RRRRzNdgRV:RFHsRRRHM5b8C0ME_kOl_C#DDR4-R2FR8IFM0RojRCsMCN
0CSR--Q5VRNs88I0H8ERR>gM2RCRC80OFRs0CNCsRIHR0CCLMNDNCRMF8Rkk0b0MRCNCLDRD#CCRO0DHFoOS
SSjzcNRR:H5VRNs88I0H8ERR>go2RCsMCN
0CSR--VRHGVRFsODNDRU4dUR(,#CCDOF0RVsR0HN#00MCRFL0RCoHMRosCHC#0s
C8SSSSs0Fk_5CMH<2R=4R''ERIC5MR)7q7)l_0b85N8HsI8-0E4FR8IFM0RRg2=2RHR#CDCjR''S;
SISSF_k0CHM52=R<R''4RCIEMIR5Ns8_CNo58I8sHE80-84RF0IMF2RgRH=RRC2RDR#C';j'
SSSS0Is_5CMH<2R= RWRCIEMIR5Ns8_CNo58I8sHE80-84RF0IMF2RgRH=R2DRC#'CRj
';SCSSMo8RCsMCNR0CzNcj;-
S-VRQR85N8HsI8R0E<g=R2FRMRHIs0CCRMDNLCsRFR0FkbRk0CLMND#CRCODC0FRDoRHOM8CCCS8
ScSz4:NRRRHV58N8s8IH0<ER=2RgRMoCC0sNCS
SSFSskC0_M25HRR<=';4'
SSSSkIF0M_C5RH2<'=R4
';SSSSI_s0CHM52=R<R;W 
SSSCRM8oCCMsCN0R4zcNS;
-t-RCsMCNR0C0REC)RqvODCD#MRN8sR0H0-#N#0C
SSSzNc.RV:RF[sRRRHM58IH0ME_kOl_C#DDR4-R2FR8IFM0RojRCsMCN
0CRRRRRRRRRRRRRRRRNs00H0LkC3R\s_NlF#VVCR0\FAVR)_qv6X4.dR.7:NRDLRCDH"#RW
";RRRRRRRRRRRRRRRRLHCoMR
RRRRRRRRRRRRRRRRRAv)q_.64X7d.R):Rq4vAnd_1nd_1nR
RRRRRRRRRRRRRRRRRRFRbsl0RN5bR7RQq=H>RMC_son5d*d[+4FR8IFM0R*dn[R2,q)77q>R=RIDF_8IN8Us5RI8FMR0FjR2,7RQA=">Rjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"q,R7A7)RR=>D_FIs8N8sR5U8MFI0jFR2R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRq hRR=>',4'R)11q>R=R''j, RWq>R=R0Is_5CMHR2,BqpiRR=>B,piRA hRR=>',4'R)11A>R=R''j, RWA>R=R''j,pRBi=AR>pRBiR,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRq7m52d4RR=>I0Fk_#LkdH.5,*d.[4+d2
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRmR7qj5d2>R=RkIF0k_L#5d.H.,d*d[+j
2,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRmR7qg5.2>R=RkIF0k_L#5d.H.,d*.[+gR2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRR7RRm.q5U=2R>FRIkL0_k.#d5dH,.+*[.,U2RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mq.R(2=I>RF_k0Ldk#.,5Hd[.*+2.(,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mq.Rn2=I>RF_k0Ldk#.,5Hd[.*+2.n,RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRq7m52.6RR=>I0Fk_#LkdH.5,*d.[6+.2
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRmR7qc5.2>R=RkIF0k_L#5d.H.,d*.[+c
2,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRmR7qd5.2>R=RkIF0k_L#5d.H.,d*.[+dR2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRR7RRm.q5.=2R>FRIkL0_k.#d5dH,.+*[.,.2RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mq.R42=I>RF_k0Ldk#.,5Hd[.*+2.4,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mq.Rj2=I>RF_k0Ldk#.,5Hd[.*+2.j,RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRq7m524gRR=>I0Fk_#LkdH.5,*d.[g+42
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRmR7qU542>R=RkIF0k_L#5d.H.,d*4[+U
2,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRmR7q(542>R=RkIF0k_L#5d.H.,d*4[+(R2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRR7RRm4q5n=2R>FRIkL0_k.#d5dH,.+*[4,n2RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mq4R62=I>RF_k0Ldk#.,5Hd[.*+246,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mq4Rc2=I>RF_k0Ldk#.,5Hd[.*+24c,RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRq7m524dRR=>I0Fk_#LkdH.5,*d.[d+42
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRmR7q.542>R=RkIF0k_L#5d.H.,d*4[+.
2,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRmR7q4542>R=RkIF0k_L#5d.H.,d*4[+4R2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRR7RRm4q5j=2R>FRIkL0_k.#d5dH,.+*[4,j2RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mqg=2R>FRIkL0_k.#d5dH,.+*[g
2,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRmR7q25URR=>I0Fk_#LkdH.5,*d.[2+U,RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRq7m5R(2=I>RF_k0Ldk#.,5Hd[.*+,(2RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mqn=2R>FRIkL0_k.#d5dH,.+*[n
2,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRmR7q256RR=>I0Fk_#LkdH.5,*d.[2+6,RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRq7m5Rc2=I>RF_k0Ldk#.,5Hd[.*+,c2RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mqd=2R>FRIkL0_k.#d5dH,.+*[d
2,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRmR7q25.RR=>I0Fk_#LkdH.5,*d.[2+.,RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRq7m5R42=I>RF_k0Ldk#.,5Hd[.*+,42RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mqj=2R>FRIkL0_k.#d5dH,.2*[,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mAdR42=s>RF_k0Ldk#.,5Hd[.*+2d4,RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRA7m52djRR=>s0Fk_#LkdH.5,*d.[j+d2R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRA7m52.gRR=>s0Fk_#LkdH.5,*d.[g+.2
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRmR7AU5.2>R=RksF0k_L#5d.H.,d*.[+UR2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRR7RRm.A5(=2R>FRskL0_k.#d5dH,.+*[.,(2
RRRRRRRRRRRRRRRRRRRRRRRRRRRR7RRm.A5n=2R>FRskL0_k.#d5dH,.+*[.,n2RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mA.R62=s>RF_k0Ldk#.,5Hd[.*+2.6,RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRA7m52.cRR=>s0Fk_#LkdH.5,*d.[c+.2R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRA7m52.dRR=>s0Fk_#LkdH.5,*d.[d+.2
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRmR7A.5.2>R=RksF0k_L#5d.H.,d*.[+.R2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRR7RRm.A54=2R>FRskL0_k.#d5dH,.+*[.,42
RRRRRRRRRRRRRRRRRRRRRRRRRRRR7RRm.A5j=2R>FRskL0_k.#d5dH,.+*[.,j2RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mA4Rg2=s>RF_k0Ldk#.,5Hd[.*+24g,RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRA7m524URR=>s0Fk_#LkdH.5,*d.[U+42R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRA7m524(RR=>s0Fk_#LkdH.5,*d.[(+42
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRmR7An542>R=RksF0k_L#5d.H.,d*4[+nR2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRR7RRm4A56=2R>FRskL0_k.#d5dH,.+*[4,62
RRRRRRRRRRRRRRRRRRRRRRRRRRRR7RRm4A5c=2R>FRskL0_k.#d5dH,.+*[4,c2RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mA4Rd2=s>RF_k0Ldk#.,5Hd[.*+24d,RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRA7m524.RR=>s0Fk_#LkdH.5,*d.[.+42R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRA7m5244RR=>s0Fk_#LkdH.5,*d.[4+42
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRmR7Aj542>R=RksF0k_L#5d.H.,d*4[+jR2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRR7RRmgA52>R=RksF0k_L#5d.H.,d*g[+2R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRA7m5RU2=s>RF_k0Ldk#.,5Hd[.*+,U2RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mA(=2R>FRskL0_k.#d5dH,.+*[(R2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRR7RRmnA52>R=RksF0k_L#5d.H.,d*n[+2R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRA7m5R62=s>RF_k0Ldk#.,5Hd[.*+,62RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mAc=2R>FRskL0_k.#d5dH,.+*[cR2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRR7RRmdA52>R=RksF0k_L#5d.H.,d*d[+2R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRA7m5R.2=s>RF_k0Ldk#.,5Hd[.*+,.2RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mA4=2R>FRskL0_k.#d5dH,.+*[4R2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRR7RRmjA52>R=RksF0k_L#5d.H.,d*,[2
RRRRRRRRRRRRRRRRRRRRRRRRRRRR7RRQRuq=H>RMC_son5d*d[+6FR8IFM0R*dn[.+d27,RQRuA=">Rjjjj"R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRu7mq25dRR=>IsbNH_0$Ldk#.,5Hc+*[dR2,7qmu5R.2=I>RbHNs0L$_k.#d5cH,*.[+2R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRu7mq254RR=>IsbNH_0$Ldk#.,5Hc+*[4R2,7qmu5Rj2=I>RbHNs0L$_k.#d5cH,*,[2
RRRRRRRRRRRRRRRRRRRRRRRRRRRR7RRm5uAd=2R>bRsN0sH$k_L#5d.H*,c[2+d,mR7u.A52>R=RNsbs$H0_#LkdH.5,[c*+,.2
RRRRRRRRRRRRRRRRRRRRRRRRRRRR7RRm5uA4=2R>bRsN0sH$k_L#5d.H*,c[2+4,mR7ujA52>R=RNsbs$H0_#LkdH.5,[c*2
2;RRRRRRRRRRRRRRRRRFRsks0_Cdo5n2*[RR<=s0Fk_#LkdH.5,*d.[I2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRsRRF_k0s5Cod[n*+R42<s=RF_k0Ldk#.,5Hd[.*+R42IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRs0Fk_osC5*dn[2+.RR<=s0Fk_#LkdH.5,*d.[2+.RCIEMsR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRksF0C_son5d*d[+2=R<RksF0k_L#5d.H.,d*d[+2ERIC5MRs0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRFRsks0_Cdo5n+*[c<2R=FRskL0_k.#d5dH,.+*[cI2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRsRRF_k0s5Cod[n*+R62<s=RF_k0Ldk#.,5Hd[.*+R62IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRs0Fk_osC5*dn[2+nRR<=s0Fk_#LkdH.5,*d.[2+nRCIEMsR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRksF0C_son5d*([+2=R<RksF0k_L#5d.H.,d*([+2ERIC5MRs0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRFRsks0_Cdo5n+*[U<2R=FRskL0_k.#d5dH,.+*[UI2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRsRRF_k0s5Cod[n*+Rg2<s=RF_k0Ldk#.,5Hd[.*+Rg2IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRs0Fk_osC5*dn[j+42=R<RksF0k_L#5d.H.,d*4[+jI2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRsRRF_k0s5Cod[n*+244RR<=s0Fk_#LkdH.5,*d.[4+42ERIC5MRs0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRFRsks0_Cdo5n+*[4R.2<s=RF_k0Ldk#.,5Hd[.*+24.RCIEMsR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRksF0C_son5d*4[+d<2R=FRskL0_k.#d5dH,.+*[4Rd2IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRs0Fk_osC5*dn[c+42=R<RksF0k_L#5d.H.,d*4[+cI2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRsRRF_k0s5Cod[n*+246RR<=s0Fk_#LkdH.5,*d.[6+42ERIC5MRs0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRFRsks0_Cdo5n+*[4Rn2<s=RF_k0Ldk#.,5Hd[.*+24nRCIEMsR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRksF0C_son5d*4[+(<2R=FRskL0_k.#d5dH,.+*[4R(2IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRs0Fk_osC5*dn[U+42=R<RksF0k_L#5d.H.,d*4[+UI2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRsRRF_k0s5Cod[n*+24gRR<=s0Fk_#LkdH.5,*d.[g+42ERIC5MRs0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRFRsks0_Cdo5n+*[.Rj2<s=RF_k0Ldk#.,5Hd[.*+2.jRCIEMsR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRksF0C_son5d*.[+4<2R=FRskL0_k.#d5dH,.+*[.R42IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRs0Fk_osC5*dn[.+.2=R<RksF0k_L#5d.H.,d*.[+.I2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRsRRF_k0s5Cod[n*+2.dRR<=s0Fk_#LkdH.5,*d.[d+.2ERIC5MRs0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRFRsks0_Cdo5n+*[.Rc2<s=RF_k0Ldk#.,5Hd[.*+2.cRCIEMsR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRksF0C_son5d*.[+6<2R=FRskL0_k.#d5dH,.+*[.R62IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRs0Fk_osC5*dn[n+.2=R<RksF0k_L#5d.H.,d*.[+nI2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRsRRF_k0s5Cod[n*+2.(RR<=s0Fk_#LkdH.5,*d.[(+.2ERIC5MRs0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRFRsks0_Cdo5n+*[.RU2<s=RF_k0Ldk#.,5Hd[.*+2.URCIEMsR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRksF0C_son5d*.[+g<2R=FRskL0_k.#d5dH,.+*[.Rg2IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRs0Fk_osC5*dn[j+d2=R<RksF0k_L#5d.H.,d*d[+jI2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRsRRF_k0s5Cod[n*+2d4RR<=s0Fk_#LkdH.5,*d.[4+d2ERIC5MRs0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRFRsks0_Cdo5n+*[dR.2<s=RbHNs0L$_k.#d5cH,*R[2IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRs0Fk_osC5*dn[d+d2=R<RNsbs$H0_#LkdH.5,[c*+R42IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRs0Fk_osC5*dn[c+d2=R<RNsbs$H0_#LkdH.5,[c*+R.2IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRs0Fk_osC5*dn[6+d2=R<RNsbs$H0_#LkdH.5,[c*+Rd2IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRR
RRRRRRRRRRRRRRRRIRRF_k0s5Cod[n*2=R<RkIF0k_L#5d.H.,d*R[2IMECRF5IkC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRI0Fk_osC5*dn[2+4RR<=I0Fk_#LkdH.5,*d.[2+4RCIEMIR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRkIF0C_son5d*.[+2=R<RkIF0k_L#5d.H.,d*.[+2ERIC5MRI0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRFRIks0_Cdo5n+*[d<2R=FRIkL0_k.#d5dH,.+*[dI2RERCM5kIF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRIRRF_k0s5Cod[n*+Rc2<I=RF_k0Ldk#.,5Hd[.*+Rc2IMECRF5IkC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRI0Fk_osC5*dn[2+6RR<=I0Fk_#LkdH.5,*d.[2+6RCIEMIR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRkIF0C_son5d*n[+2=R<RkIF0k_L#5d.H.,d*n[+2ERIC5MRI0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRFRIks0_Cdo5n+*[(<2R=FRIkL0_k.#d5dH,.+*[(I2RERCM5kIF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRIRRF_k0s5Cod[n*+RU2<I=RF_k0Ldk#.,5Hd[.*+RU2IMECRF5IkC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRI0Fk_osC5*dn[2+gRR<=I0Fk_#LkdH.5,*d.[2+gRCIEMIR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRkIF0C_son5d*4[+j<2R=FRIkL0_k.#d5dH,.+*[4Rj2IMECRF5IkC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRI0Fk_osC5*dn[4+42=R<RkIF0k_L#5d.H.,d*4[+4I2RERCM5kIF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRIRRF_k0s5Cod[n*+24.RR<=I0Fk_#LkdH.5,*d.[.+42ERIC5MRI0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRFRIks0_Cdo5n+*[4Rd2<I=RF_k0Ldk#.,5Hd[.*+24dRCIEMIR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRkIF0C_son5d*4[+c<2R=FRIkL0_k.#d5dH,.+*[4Rc2IMECRF5IkC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRI0Fk_osC5*dn[6+42=R<RkIF0k_L#5d.H.,d*4[+6I2RERCM5kIF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRIRRF_k0s5Cod[n*+24nRR<=I0Fk_#LkdH.5,*d.[n+42ERIC5MRI0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRFRIks0_Cdo5n+*[4R(2<I=RF_k0Ldk#.,5Hd[.*+24(RCIEMIR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRkIF0C_son5d*4[+U<2R=FRIkL0_k.#d5dH,.+*[4RU2IMECRF5IkC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRI0Fk_osC5*dn[g+42=R<RkIF0k_L#5d.H.,d*4[+gI2RERCM5kIF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRIRRF_k0s5Cod[n*+2.jRR<=I0Fk_#LkdH.5,*d.[j+.2ERIC5MRI0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRFRIks0_Cdo5n+*[.R42<I=RF_k0Ldk#.,5Hd[.*+2.4RCIEMIR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRkIF0C_son5d*.[+.<2R=FRIkL0_k.#d5dH,.+*[.R.2IMECRF5IkC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRI0Fk_osC5*dn[d+.2=R<RkIF0k_L#5d.H.,d*.[+dI2RERCM5kIF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRIRRF_k0s5Cod[n*+2.cRR<=I0Fk_#LkdH.5,*d.[c+.2ERIC5MRI0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRFRIks0_Cdo5n+*[.R62<I=RF_k0Ldk#.,5Hd[.*+2.6RCIEMIR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRkIF0C_son5d*.[+n<2R=FRIkL0_k.#d5dH,.+*[.Rn2IMECRF5IkC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRI0Fk_osC5*dn[(+.2=R<RkIF0k_L#5d.H.,d*.[+(I2RERCM5kIF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRIRRF_k0s5Cod[n*+2.URR<=I0Fk_#LkdH.5,*d.[U+.2ERIC5MRI0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRFRIks0_Cdo5n+*[.Rg2<I=RF_k0Ldk#.,5Hd[.*+2.gRCIEMIR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRkIF0C_son5d*d[+j<2R=FRIkL0_k.#d5dH,.+*[dRj2IMECRF5IkC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRI0Fk_osC5*dn[4+d2=R<RkIF0k_L#5d.H.,d*d[+4I2RERCM5kIF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRIRRF_k0s5Cod[n*+2d.RR<=IsbNH_0$Ldk#.,5Hc2*[RCIEMIR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRkIF0C_son5d*d[+d<2R=bRIN0sH$k_L#5d.H*,c[2+4RCIEMIR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRkIF0C_son5d*d[+c<2R=bRIN0sH$k_L#5d.H*,c[2+.RCIEMIR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRkIF0C_son5d*d[+6<2R=bRIN0sH$k_L#5d.H*,c[2+dRCIEMIR5F_k0CHM52RR='24'R#CDCZR''
;
SCSSMo8RCsMCNR0CzNc.;S
SCRM8oCCMsCN0RgzdNS;
CRM8oCCMsCN0RUzdNR;
R8CMRMoCC0sNCcRzd
;
RcRzcRR:H5VRMRF0s8N8sC_soo2RCsMCNR0C-o-RCsMCNR0C#CCDOs0RNRl
R-RR-VRQR8N8s8IH0<ERRN6R#o#HMjR''FR0RkkM#RC8L#H0
RRRRRzjRH:RVNR58I8sHE80R4=R2CRoMNCs0RC
RRRRRDRRFsI_Ns88_<#R=jR"jjjj"RR&s_N8s_Co#25j;R
RRRRRRFRDIN_I8_8s#=R<Rj"jj"jjRI&RNs8_C#o_5;j2
RRRR8CMRMoCC0sNCjRz;R
RR4RzRRR:H5VRNs88I0H8ERR=.o2RCsMCN
0CRRRRRRRRD_FIs8N8sR_#<"=Rjjjj"RR&s_N8s_Co#R548MFI0jFR2R;
RRRRRDRRFII_Ns88_<#R=jR"j"jjRI&RNs8_C#o_584RF0IMF2Rj;R
RRMRC8CRoMNCs0zCR4R;
RzRR.:RRRRHV58N8s8IH0=ERRRd2oCCMsCN0
RRRRRRRRIDF_8sN8#s_RR<="jjj"RR&s_N8s_Co#R5.8MFI0jFR2R;
RRRRRDRRFII_Ns88_<#R=jR"jRj"&NRI8C_so5_#.FR8IFM0R;j2
RRRR8CMRMoCC0sNC.Rz;R
RRdRzRRR:H5VRNs88I0H8ERR=co2RCsMCN
0CRRRRRRRRD_FIs8N8sR_#<"=RjRj"&NRs8C_so5_#dFR8IFM0R;j2
RRRRRRRRIDF_8IN8#s_RR<=""jjRI&RNs8_C#o_58dRF0IMF2Rj;R
RRMRC8CRoMNCs0zCRdS;
z:cSRRHV58N8s8IH0=ERRR62oCCMsCN0
DSSFsI_Ns88_<#R=jR''RR&s_N8s_Co#R5c8MFI0jFR2S;
SIDF_8IN8#s_RR<='Rj'&NRI8C_so5_#cFR8IFM0R;j2
MSC8CRoMNCs0zCRcR;
RzRR6:RRRRHV58N8s8IH0>ERRR62oCCMsCN0
RRRRRRRRIDF_8sN8#s_RR<=s_N8s_Co#R568MFI0jFR2R;
RRRRRDRRFII_Ns88_<#R=NRI8C_so5_#6FR8IFM0R;j2
RRRR8CMRMoCC0sNC6Rz;R

R-RR-VRQRH58MC_sos2RC#oH0RCs7RQhkM#HopRBiR
RRnRzRRR:H5VR8_HMs2CoRMoCC0sNCR
RRRRRRsRbF#OC#BR5pRi,72QhRoLCHRM
RRRRRRRRRHRRVBR5p=iRR''4R8NMRiBp'CCPMR020MEC
RRRRRRRRRRRRRRRR_HMs_Co#=R<Rh7Q;R
RRRRRRRRRRMRC8VRH;R
RRRRRRMRC8sRbF#OC#R;
RCRRMo8RCsMCNR0Cz
n;RRRRzR(R:VRHRF5M0HR8MC_soo2RCsMCN
0CRRRRRRRRRRRRHsM_C#o_RR<=7;Qh
RRRR8CMRMoCC0sNC(Rz;R

R-RR-VRQR85sF_k0s2CoRosCHC#0smR7zkaR#oHMRpmBiR
RRURzs:RRRRHV5Fs8ks0_CRo2oCCMsCN0
RRRRRRRRFbsO#C#R_5)miBp,FRsks0_C#o_2CRLo
HMRRRRRRRRRRRRH5VR)B_mp=iRR''4R8NMRm)_B'piCMPC002RE
CMRRRRRRRRRRRRRRRR)m_7z<aR=FRsks0_C#o_;R
RRRRRRRRRRMRC8VRH;R
RRRRRRMRC8sRbF#OC#R;
RCRRMo8RCsMCNR0Cz;Us
RRRRszgRRR:H5VRMRF0sk8F0C_soo2RCsMCN
0CRRRRRRRRRRRR)m_7z<aR=FRsks0_C#o_;R
RRMRC8CRoMNCs0zCRg
s;
USzI:RRRRHV5FI8ks0_CRo2oCCMsCN0
RRRRRRRRFbsO#C#R_5WmiBp,FRIks0_C#o_2CRLo
HMRRRRRRRRRRRRH5VRWB_mp=iRR''4R8NMRmW_B'piCMPC002RE
CMRRRRRRRRRRRRRRRRWm_7z<aR=FRIks0_C#o_;R
RRRRRRRRRRMRC8VRH;R
RRRRRRMRC8sRbF#OC#R;
RCRRMo8RCsMCNR0Cz;UI
RRRRIzgRRR:H5VRMRF0Ik8F0C_soo2RCsMCN
0CRRRRRRRRRRRRWm_7z<aR=FRIks0_C#o_;R
RRMRC8CRoMNCs0zCRg
I;
RRRRR--Q5VRs8N8sC_sos2RC#oH0RCsq)77RHk#MBoRpRi
RzRR4RjR:VRHRN5s8_8ss2CoRMoCC0sNCR
RRRRRRsRbF#OC#)R5_pmBi),Rq)772CRLo
HMRRRRRRRRRRRRH5VR)B_mp=iRR''4R8NMRm)_B'piCMPC002RE
CMRRRRRRRRRRRRRRRRs_N8s_Co#=R<R7)q7N)58I8sHE80-84RF0IMF2Rj;R
RRRRRRRRRRMRC8VRH;R
RRRRRRMRC8sRbF#OC#R;
RCRRMo8RCsMCNR0Cz;4j
RRRR4z4RH:RVMR5Fs0RNs88_osC2CRoMNCs0RC
RRRRRRRRRsRRNs8_C#o_RR<=)7q7)R;
RCRRMo8RCsMCNR0Cz;44
R
RR-R-RRQV58IN8ss_CRo2sHCo#s0CR7q7)#RkHRMoB
piRRRRzR4.RH:RVIR5Ns88_osC2CRoMNCs0RC
RRRRRbRRsCFO#5#RB,piR7Wq7R)2LHCoMR
RRRRRRRRRRVRHRp5BiRR='R4'NRM8B'piCMPC002RE
CMRRRRRRRRRRRRRRRRI_N8s_Co#=R<R7Wq7N)58I8sHE80-84RF0IMF2Rj;R
RRRRRRRRRRMRC8VRH;R
RRRRRRMRC8sRbF#OC#R;
RCRRMo8RCsMCNR0Cz;4.
RRRRdz4RH:RVMR5FI0RNs88_osC2CRoMNCs0RC
RRRRRRRRRIRRNs8_C#o_RR<=W7q7)R;
RCRRMo8RCsMCNR0Cz;4d
RRRRRRRRR
RR-R-RMtCC0sNCER0CqR)vCRODRD#NRM8#CCDOD0RFOoH
RRRRcz4RV:RFHsRRRHM5lMk_DOCDc_nR4-R2FR8IFM0RojRCsMCN
0CRRRR-Q-RVNR58I8sHE80R6>R2CRMC08RFsROCCN0RHIs0CCRMDNLCMRN8kRF00bkRNCMLRDC#CCDOD0RFOoH
RRRRRRRR6z4RH:RVNR58I8sHE80Rn>R2CRoMNCs0RC
RRRRRRRRRRRRRsRRF_k0C#M_5RH2<'=R4I'RERCM58sN_osC_N#58I8sHE80-84RF0IMF2RnRH=R2DRC#'CRj
';SSSSI0Fk__CM#25HRR<='R4'IMECRN5I8C_so5_#Ns88I0H8ER-48MFI0nFR2RR=HC2RDR#C';j'
RRRRRRRRRRRRRRRR0Is__CM#25HRR<=WI RERCM58IN_osC_N#58I8sHE80-84RF0IMF2RnRH=R2DRC#'CRj
';RRRRRRRRCRM8oCCMsCN0R6z4;R
RR-R-RRQV58N8s8IH0<ER=2R6RRMFI0sHCMRCNCLDRRFsFbk0kC0RMDNLCCR#D0CORoDFHMORCCC88R
RRRRRR4RznRR:H5VRNs88I0H8E=R<RRn2oCCMsCN0
RRRRRRRRRRRRRRRRksF0M_C_H#52=R<R''4;S
SSFSIkC0_M5_#H<2R=4R''R;
RRRRRRRRRRRRRIRRsC0_M5_#H<2R= RW;R
RRRRRRMRC8CRoMNCs0zCR4
n;RRRR-t-RCsMCNR0C0REC)RqvODCD#MRN8sR0H0-#N#0C
RRRRRRRR(z4RV:RF[sRRRHM58IH0-ERRR428MFI0jFRRMoCC0sNCR
RRRRRRRRRR0RN0LsHkR0C\N3slV_FV0#C\VRFRqz)vRnc:NRDLRCDH"#R1"7aRH&RMo0CCHs'lCNo58IH0RE2&7R""RR&HCM0o'CsHolNC*5HnRc2&WR""RR&HCM0o'CsHolNC25[R"&R &"RR0HMCsoC'NHlooC5CC0_M88_CEb05+5H4n2*c8,RCEb02&2RR""XRH&RMo0CCHs'lCNo54[+2R;
RRRRRRRRRLRRCMoH
RRRRRRRRRRRRqz)vRnc:)RXqcvnXR47
RRRRRRRRRRRRRRRRsbF0NRlb7R5RR=>HsM_C#o_5,[2RRqj=D>RFII_Ns88_j#52q,R4>R=RIDF_8IN8#s_5,42RRq.=D>RFII_Ns88_.#52R,
RRRRRRRRRRRRRRRRRRRRRRRRRRqd=D>RFII_Ns88_d#52q,Rc>R=RIDF_8IN8#s_5,c2RRq6=D>RFII_Ns88_6#52
,RSSSSSRSR7qu)j>R=RIDF_8sN8#s_5,j2R)7uq=4R>FRDIN_s8_8s#254,uR7)Rq.=D>RFsI_Ns88_.#52S,
SSSSS7RRud)qRR=>D_FIs8N8s5_#dR2,7qu)c>R=RIDF_8sN8#s_5,c2R)7uq=6R>FRDIN_s8_8s#256,SR
SSSSSWRR >R=R0Is__CM#25H,BRWp=iR>pRBi7,Ru=mR>FRskL0_kn#_cH#5,,[2Rm1uRR=>I0Fk_#Lk_#nc5[H,2
2;RRRRRRRRRRRRRRRRs0Fk_osC_[#52=R<RksF0k_L#c_n#,5H[I2RERCM5ksF0M_C_H#52RR='24'R#CDCZR''S;
SISSF_k0s_Co#25[RR<=I0Fk_#Lk_#nc5[H,2ERIC5MRI0Fk__CM#25HR'=R4R'2CCD#R''Z;R
RRRRRRMRC8CRoMNCs0zCR4
(;RRRRR8CMRMoCC0sNC4RzcR;RRRRRRRRRRRR
RRRRRR
RR-R-RMtCC0sNCRRNdI.RFRs88bCCRv)qRDOCDVRHRbNbssFbHCN0RRRRRRRRRRRRR
RRRRRRzR4U:VRHRk5MlC_ODdD_.RR=4o2RCsMCN
0CRRRR-Q-RVNR58I8sHE80R(>R2CRMC08RFsROCCN0RHIs0CCRMDNLCMRN8kRF00bkRNCMLRDC#CCDOD0RFOoH
RRRRRRRRgz4NRR:H5VRNs88I0H8ERR>no2RCsMCN
0CRRRRRRRRRRRRRRRRs0Fk__CMd<.R=4R''ERIC5MR58sN_osC_N#58I8sHE80-84RF0IMF2RnRM=RkOl_C_DDnRc2NRM858sN_osC_6#52RR='2j'2DRC#'CRj
';SSSSI0Fk__CMd<.R=4R''ERIC5MR58IN_osC_N#58I8sHE80-84RF0IMF2RnRM=RkOl_C_DDnRc2NRM858IN_osC_6#52RR='2j'2DRC#'CRj
';RRRRRRRRRRRRRRRRI_s0CdM_.=R<RRW IMECRI55Ns8_C#o_58N8s8IH04E-RI8FMR0Fn=2RRlMk_DOCDc_n2MRN8IR5Ns8_C#o_5R62=jR''R22CCD#R''j;R
RRRRRRMRC8CRoMNCs0zCR4;gN
RRRRRRRRgz4LRR:H5VRNs88I0H8ERR=nMRN8kRMlC_ODnD_cRR=jo2RCsMCN
0CRRRRRRRRRRRRRRRRs0Fk__CMd<.R=4R''ERIC5MR58sN_osC_6#52RR='2j'2DRC#'CRj
';SSSSI0Fk__CMd<.R=4R''ERIC5MR58IN_osC_6#52RR='2j'2DRC#'CRj
';RRRRRRRRRRRRRRRRI_s0CdM_.=R<RRW IMECRI55Ns8_C#o_5R62=jR''R22CCD#R''j;R
RRRRRRMRC8CRoMNCs0zCR4;gLRRRR-Q-RVNR58I8sHE80RR<=6M2RFsRIHR0CCLMNDFCRskRF00bkRNCMLRDC#CCDOD0RFOoHRCMC8
C8RRRRRRRRzR.j:VRHR85N8HsI8R0E<6=R2CRoMNCs0RC
RRRRRRRRRRRRRsRRF_k0CdM_.=R<R''4;S
SSFSIkC0_M._dRR<=';4'
RRRRRRRRRRRRRRRR0Is__CMd<.R= RW;R
RRRRRRMRC8CRoMNCs0zCR.
j;RRRR-t-RCsMCNR0C0REC)RqvODCDR8NMRH0s-N#00RC
RRRRRzRR.:4RRsVFRH[RMIR5HE80R4-R2FR8IFM0RojRCsMCN
0CRRRRRRRRRRRRNs00H0LkC3R\s_NlF#VVCR0\FzVR)dqv.RR:DCNLD#RHR7"1a&"RR0HMCsoC'NHloIC5HE802RR&"R7"&MRH0CCosl'HN5oCM_klODCD_*ncnRc2&WR""RR&HCM0o'CsHolNC25[R"&R &"RR0HMCsoC'NHlooC5CC0_M88_CEb05lMk_DOCDc_n*Rnc+.Rd,CR8b20E2RR&"RX"&MRH0CCosl'HN5oC[2+4;R
RRRRRRRRRRCRLo
HMRRRRRRRRRRRRzv)qd:.RRqX)vXd.4
7RRRRRRRRRRRRRRRRRb0FsRblNRR57=H>RMC_so5_#[R2,q=jR>FRDIN_I8_8s#25j,4RqRR=>D_FII8N8s5_#4R2,q=.R>FRDIN_I8_8s#25.,R
RRRRRRRRRRRRRRRRRRRRRRRRRq=dR>FRDIN_I8_8s#25d,cRqRR=>D_FII8N8s5_#cR2,
SSSSRSSR)7uq=jR>FRDIN_s8_8s#25j,uR7)Rq4=D>RFsI_Ns88_4#527,Ru.)qRR=>D_FIs8N8s5_#.
2,SSSSSRSR7qu)d>R=RIDF_8sN8#s_5,d2R)7uq=cR>FRDIN_s8_8s#25c,SR
SSSSSWRR >R=R0Is__CMdR.,WiBpRR=>B,piRm7uRR=>s0Fk_#Lk_#d.5lMk_DOCD._d,,[2Rm1uRR=>I0Fk_#Lk_#d.5lMk_DOCD._d,2[2;R
RRRRRRRRRRRRRRFRsks0_C#o_5R[2<s=RF_k0L_k#d5.#M_klODCD_,d.[I2RERCM5ksF0M_C_Rd.=4R''C2RDR#C';Z'
SSSSkIF0C_so5_#[<2R=FRIkL0_kd#_.M#5kOl_C_DDd[.,2ERIC5MRI0Fk__CMd=.RR''42DRC#'CRZ
';RRRRRRRRR8CMRMoCC0sNC.Rz4R;
RRRRCRM8oCCMsCN0RUz4;RRRRRRRR
RR
RRRRR--tCCMsCN0R4NRnFRIs88RCRCb)RqvODCDRRHVNsbbFHbsNR0CRRRRRRRRRRRRRRR
RzRR.:.RRRHV5lMk_DOCDn_4R4=R2CRoMNCs0RC
R-RR-VRQR85N8HsI8R0E>2R6RCMC8FR0RCOsNR0CI0sHCMRCNCLDR8NMR0FkbRk0CLMND#CRCODC0FRDo
HORRRRRRRRzN.dRH:RVNR58I8sHE80Rn>RR8NMRlMk_DOCD._dR4=R2CRoMNCs0RC
RRRRRRRRRRRRRsRRF_k0C4M_n=R<R''4RCIEM5R5s_N8s_Co#85N8HsI8-0E4FR8IFM0RRn2=kRMlC_ODnD_cN2RM58Rs_N8s_Co#256R'=R4R'2NRM858sN_osC_c#52RR='2j'2DRC#'CRj
';SSSSI0Fk__CM4<nR=4R''ERIC5MR58IN_osC_N#58I8sHE80-84RF0IMF2RnRM=RkOl_C_DDnRc2NRM858IN_osC_6#52RR='24'R8NMRN5I8C_so5_#c=2RR''j2C2RDR#C';j'
RRRRRRRRRRRRRRRR0Is__CM4<nR= RWRCIEM5R5I_N8s_Co#85N8HsI8-0E4FR8IFM0RRn2=kRMlC_ODnD_cN2RM58RI_N8s_Co#256R'=R4R'2NRM858IN_osC_c#52RR='2j'2DRC#'CRj
';RRRRRRRRCRM8oCCMsCN0Rdz.NR;
RRRRRzRR.RdL:VRHR85N8HsI8R0E>RRnNRM8M_klODCD_Rd./4=R2CRoMNCs0RC
RRRRRRRRRRRRRsRRF_k0C4M_n=R<R''4RCIEM5R5s_N8s_Co#85N8HsI8-0E4FR8IFM0RRn2=kRMlC_ODnD_cN2RM58Rs_N8s_Co#256R'=RjR'2NRM858sN_osC_c#52RR='2j'2DRC#'CRj
';SSSSI0Fk__CM4<nR=4R''ERIC5MR58IN_osC_N#58I8sHE80-84RF0IMF2RnRM=RkOl_C_DDnRc2NRM858IN_osC_6#52RR='2j'R8NMRN5I8C_so5_#c=2RR''j2C2RDR#C';j'
RRRRRRRRRRRRRRRR0Is__CM4<nR= RWRCIEM5R5I_N8s_Co#85N8HsI8-0E4FR8IFM0RRn2=kRMlC_ODnD_cN2RM58RI_N8s_Co#256R'=RjR'2NRM858IN_osC_c#52RR='2j'2DRC#'CRj
';RRRRRRRRCRM8oCCMsCN0Rdz.LR;
RRRRRzRR.RdO:VRHR85N8HsI8R0E=RRnNRM8M_klODCD_Rd.=2R4RMoCC0sNCR
RRRRRRRRRRRRRRFRskC0_Mn_4RR<='R4'IMECRs55Ns8_C#o_5R62=4R''N2RM58Rs_N8s_Co#25cR'=Rj2'2R#CDCjR''S;
SISSF_k0C4M_n=R<R''4RCIEM5R5I_N8s_Co#256R'=R4R'2NRM858IN_osC_c#52RR='2j'2DRC#'CRj
';RRRRRRRRRRRRRRRRI_s0C4M_n=R<RRW IMECRI55Ns8_C#o_5R62=4R''N2RM58RI_N8s_Co#25cR'=Rj2'2R#CDCjR''R;
RRRRRCRRMo8RCsMCNR0CzO.d;R
RRRRRR.Rzd:8RRRHV58N8s8IH0=ERRN6RMM8RkOl_C_DDd/.R=2R4RMoCC0sNCR
RRRRRRRRRRRRRRFRskC0_Mn_4RR<='R4'IMECRs55Ns8_C#o_58N8s8IH04E-RI8FMR0Fc=2RRlMk_DOCD._d2C2RDR#C';j'
SSSSkIF0M_C_R4n<'=R4I'RERCM5N5I8C_so5_#Ns88I0H8ER-48MFI0cFR2RR=M_klODCD_2d.2DRC#'CRj
';RRRRRRRRRRRRRRRRI_s0C4M_n=R<RRW IMECRI55Ns8_C#o_58N8s8IH04E-RI8FMR0Fc=2RRlMk_DOCD._d2C2RDR#C';j'
RRRRRRRR8CMRMoCC0sNC.RzdR8;R-RR-VRQR85N8HsI8R0E<6=R2FRMRHIs0CCRMDNLCsRFR0FkbRk0CLMND#CRCODC0FRDoRHOM8CCCR8
RRRRRzRR.:cRRRHV58N8s8IH0<ER=2RcRMoCC0sNCR
RRRRRRRRRRRRRRFRskC0_Mn_4RR<=';4'
SSSSkIF0M_C_R4n<'=R4
';RRRRRRRRRRRRRRRRI_s0C4M_n=R<R;W 
RRRRRRRR8CMRMoCC0sNC.RzcR;
R-RR-CRtMNCs00CRE)CRqOvRCRDDNRM80-sH#00NCR
RRRRRR.Rz6RR:VRFs[MRHRH5I8R0E-2R4RI8FMR0FjCRoMNCs0RC
RRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)Rzqnv4RD:RNDLCRRH#"a17"RR&HCM0o'CsHolNCH5I820ER"&R7&"RR0HMCsoC'NHloMC5kOl_C_DDnnc*cRR+M_klODCD_*d.dR.2&WR""RR&HCM0o'CsHolNC25[R"&R &"RR0HMCsoC'NHlooC5CC0_M88_CEb05lMk_DOCDc_n*Rnc+kRMlC_ODdD_..*dR4+Rn8,RCEb02&2RR""XRH&RMo0CCHs'lCNo54[+2R;
RRRRRRRRRLRRCMoH
RRRRRRRRRRRRqz)vR4n:qR)vX4n4
7RRRRRRRRRRRRRRRRRb0FsRblNRR57=H>RMC_so5_#[R2,q=jR>FRDIN_I8_8s#25j,4RqRR=>D_FII8N8s5_#4R2,q=.R>FRDIN_I8_8s#25.,R
RRRRRRRRRRRRRRRRRRRRRRRRRq=dR>FRDIN_I8_8s#25d,uR7)Rqj=D>RFsI_Ns88_j#527,Ru4)qRR=>D_FIs8N8s5_#4R2,7qu).>R=RIDF_8sN8#s_5,.2
SSSSRSSR)7uq=dR>FRDIN_s8_8s#25d, RWRR=>I_s0C4M_nW,RBRpi=B>RpRi,7Rum=s>RF_k0L_k#45n#M_klODCD_,4n[R2,1Rum=I>RF_k0L_k#45n#M_klODCD_,4n[;22
RRRRRRRRRRRRRRRRksF0C_so5_#[<2R=FRskL0_k4#_nM#5kOl_C_DD4[n,2ERIC5MRs0Fk__CM4=nRR''42DRC#'CRZ
';SSSSI0Fk_osC_[#52=R<RkIF0k_L#n_4#k5MlC_OD4D_n2,[RCIEMIR5F_k0C4M_nRR='24'R#CDCZR''R;
RRRRRCRRMo8RCsMCNR0Cz;.6
RRRR8CMRMoCC0sNC.Rz.R;RRRR
R8CMRMoCC0sNCcRzcC;
MN8RsHOE00COkRsCLODF	N_sl
;
------------------------MsF_IE_OC-O	---------------------
--
ONsECH0Os0kCFRM__sIOOEC	VRFRv)q_u)W_H)R#F
OlMbFCRM0Xv)qd4.X7RRRb0FsRR5
RRRRR7RRuRmRRF:Rk#0R0k8_DHFoOR;RRRRRRRR
RRRRR1RRuRmRRF:Rk#0R0k8_DHFoO
;
RRRRRRRRqRjRRRR:H#MR0k8_DHFoOR;
RRRRRqRR4RRRRH:RM0R#8D_kFOoH;R
RRRRRR.RqRRRR:MRHR8#0_FkDo;HO
RRRRRRRRRqdR:RRRRHM#_08koDFH
O;RRRRRRRRqRcRRRR:H#MR0k8_DHFoOR;
RRRRR7RRRRRRRH:RM0R#8D_kFOoH;R
RRRRRRuR7)Rqj:MRHR8#0_FkDo;HO
RRRRRRRR)7uq:4RRRHM#_08koDFH
O;RRRRRRRR7qu).RR:H#MR0k8_DHFoOR;
RRRRR7RRud)qRH:RM0R#8D_kFOoH;R
RRRRRRuR7)Rqc:MRHR8#0_FkDo;HO
RRRRRRRRpWBi:RRRRHM#_08koDFHRO;RRRRR
RRRRRRRRRRWR RRRR:H#MR0k8_DHFoOR
RRRRRRR2;RM
C8FROlMbFC;M0
lOFbCFMMX0R)nqvc7X4RbRRFRs05R
RRRRRRuR7mRRR:kRF00R#8D_kFOoH;RRRRRRRRR
RRRRRRuR1mRRR:kRF00R#8D_kFOoH;R

RRRRRqRRjRRRRH:RM0R#8D_kFOoH;R
RRRRRR4RqRRRR:MRHR8#0_FkDo;HO
RRRRRRRRRq.R:RRRRHM#_08koDFH
O;RRRRRRRRqRdRRRR:H#MR0k8_DHFoOR;
RRRRRqRRcRRRRH:RM0R#8D_kFOoH;R
RRRRRR6RqRRRR:MRHR8#0_FkDo;HO
RRRRRRRRR7RR:RRRRHM#_08koDFH
O;RRRRRRRR7qu)jRR:H#MR0k8_DHFoOR;
RRRRR7RRu4)qRH:RM0R#8D_kFOoH;R
RRRRRRuR7)Rq.:MRHR8#0_FkDo;HO
RRRRRRRR)7uq:dRRRHM#_08koDFH
O;RRRRRRRR7qu)cRR:H#MR0k8_DHFoOR;
RRRRR7RRu6)qRH:RM0R#8D_kFOoH;R
RRRRRRBRWpRiR:MRHR8#0_FkDo;HORRRRRRRR
RRRRRRRRRW R:RRRRHM#_08koDFHRO
RRRRR;R2RCR
MO8RFFlbM0CM;k
VMHO0FVMRk_MOH0MH5:LRRFLFDMCN2CRs0MksRs#0HRMoHL#
CMoH
HRRVLR52ER0CRM
RsRRCs0kM"5"2R;
R#CDCR
RRCRs0Mks5F"BkRD8MRF0HDlbCMlC0DRAFRO	)3qvRRQ#0RECs8CNR8N8s#C#RosCHC#0sRC8kM#HoER0CNR#lOCRD	FORRN#0REC)?qv"
2;RMRC8VRH;M
C8kRVMHO_M;H0
MVkOF0HMCRo0M_C8C_8b50E#CHxRH:RMo0CC;sRRb8C0:ERR0HMCsoC2CRs0MksR0HMCsoCR
H#PHNsNCLDRMlH_x#HCRR:HCM0oRCs:j=R;C
Lo
HMRHRlMH_#x:CR=CR8b;0E
HRRV#R5HRxC<CR8b20ERC0EMR
RRHRlMH_#x:CR=HR#x
C;RMRC8VRH;R
RskC0slMRH#M_H;xC
8CMR0oC_8CM_b8C0
E;Ns00H0LkCCRoMNCs0_FssFCbs:0RRs#0H;Mo
0N0skHL0oCRCsMCNs0F_bsCFRs0FMVRFI_s_COEO:	RRONsECH0Os0kC#RHRMVkOM_HHs05Ns88_osC2-;
-CRLoRHMLODF	NRsllRHblDCCNM00MHFRo#HM#ND
b0$CMRH0s_NsRN$HN#Rs$sNRR5j06FR2VRFR0HMCsoC;F
OMN#0MI0RHE80_sNsN:$RR0HM_sNsN:$R=4R5,,R.RRc,g4,RUd,Rn
2;O#FM00NMRb8C0NE_s$sNRH:RMN0_s$sNRR:=5d4nURc,U.4g,jRcgRn,.Ujc,jR4.Rc,624.;F
OMN#0M80RH.PdRH:RMo0CC:sR=IR5HE80-/42d
n;O#FM00NMRP8H4:nRR0HMCsoCRR:=58IH04E-2U/4;F
OMN#0M80RHRPU:MRH0CCos=R:RH5I8-0E4g2/;F
OMN#0M80RHRPc:MRH0CCos=R:RH5I8-0E4c2/;F
OMN#0M80RHRP.:MRH0CCos=R:RH5I8-0E4.2/;F
OMN#0M80RHRP4:MRH0CCos=R:RH5I8-0E442/;O

F0M#NRM0LDFF4RR:LDFFCRNM:5=R84HPRj>R2O;
F0M#NRM0LDFF.RR:LDFFCRNM:5=R8.HPRj>R2O;
F0M#NRM0LDFFcRR:LDFFCRNM:5=R8cHPRj>R2O;
F0M#NRM0LDFFURR:LDFFCRNM:5=R8UHPRj>R2O;
F0M#NRM0LDFF4:nRRFLFDMCNRR:=5P8H4>nRR;j2
MOF#M0N0FRLF.DdRL:RFCFDN:MR=8R5H.PdRj>R2
;
O#FM00NMRP8H4UndcRR:HCM0oRCs:5=R80CbE2-4/d4nU
c;O#FM00NMRP8HU.4gRH:RMo0CC:sR=8R5CEb0-/42U.4g;F
OMN#0M80RHjPcg:nRR0HMCsoCRR:=5b8C04E-2j/cg
n;O#FM00NMRP8H.UjcRH:RMo0CC:sR=8R5CEb0-/42.Ujc;F
OMN#0M80RHjP4.:cRR0HMCsoCRR:=5b8C04E-2j/4.
c;O#FM00NMRP8H6R4.:MRH0CCos=R:RC58b-0E462/4
.;
MOF#M0N0FRLF4D6.RR:LDFFCRNM:5=R86HP4>.RR;j2
MOF#M0N0FRLFjD4.:cRRFLFDMCNRR:=5P8H4cj.Rj>R2O;
F0M#NRM0LDFF.UjcRL:RFCFDN:MR=8R5HjP.c>URR;j2
MOF#M0N0FRLFjDcg:nRRFLFDMCNRR:=5P8HcnjgRj>R2O;
F0M#NRM0LDFFU.4gRL:RFCFDN:MR=8R5H4PUg>.RR;j2
MOF#M0N0FRLFnD4dRUc:FRLFNDCM=R:RH58Pd4nU>cRR;j2
F
OMN#0M#0RkIl_HE80RH:RMo0CC:sR=mRAmqp hF'b#F5LF2D4RA+Rm mpqbh'FL#5F.FD2RR+Apmm 'qhb5F#LDFFc+2RRmAmph q'#bF5FLFDRU2+mRAmqp hF'b#F5LFnD42O;
F0M#NRM0#_kl80CbERR:HCM0oRCs:6=RR5-RApmm 'qhb5F#LDFF624.RA+Rm mpqbh'FL#5F4FDj2.cRA+Rm mpqbh'FL#5F.FDj2cURA+Rm mpqbh'FL#5FcFDj2gnRA+Rm mpqbh'FL#5FUFD42g.2
;
O#FM00NMROI_EOFHCH_I8R0E:MRH0CCos=R:R8IH0NE_s$sN5l#k_8IH0;E2
MOF#M0N0_RIOHEFO8C_CEb0RH:RMo0CC:sR=CR8b_0ENNss$k5#lH_I820E;F
OMN#0M80R_FOEH_OCI0H8ERR:HCM0oRCs:I=RHE80_sNsN#$5k8l_CEb02O;
F0M#NRM08E_OFCHO_b8C0:ERR0HMCsoCRR:=80CbEs_Ns5N$#_kl80CbE
2;
MOF#M0N0_RII0H8Ek_MlC_ODRD#:MRH0CCos=R:RH5I8-0E4I2/_FOEH_OCI0H8ERR+4O;
F0M#NRM0IC_8b_0EM_klODCD#RR:HCM0oRCs:5=R80CbE2-4/OI_EOFHCC_8bR0E+;R4
F
OMN#0M80R_8IH0ME_kOl_C#DDRH:RMo0CC:sR=IR5HE80-/428E_OFCHO_8IH0+ERR
4;O#FM00NMR88_CEb0_lMk_DOCD:#RR0HMCsoCRR:=5b8C04E-2_/8OHEFO8C_CEb0R4+R;O

F0M#NRM0IH_#x:CRR0HMCsoCRR:=IH_I8_0EM_klODCD#RR*IC_8b_0EM_klODCD#O;
F0M#NRM08H_#x:CRR0HMCsoCRR:=8H_I8_0EM_klODCD#RR*8C_8b_0EM_klODCD#
;
O#FM00NMRFLFDR_8:FRLFNDCM=R:R_58#CHxRI-R_x#HC=R<R;j2
MOF#M0N0FRLFID_RL:RFCFDN:MR=FRM0F5LF8D_2
;
O#FM00NMRFOEH_OCI0H8ERR:HCM0oRCs:5=RApmm 'qhb5F#LDFF_R82*_R8OHEFOIC_HE802RR+5mAmph q'#bF5FLFD2_IRI*R_FOEH_OCI0H8E
2;O#FM00NMRFOEH_OC80CbERR:HCM0oRCs:5=RApmm 'qhb5F#LDFF_R82*_R8OHEFO8C_CEb02RR+5mAmph q'#bF5FLFD2_IRI*R_FOEH_OC80CbE
2;O#FM00NMR8IH0ME_kOl_C#DDRH:RMo0CC:sR=AR5m mpqbh'FL#5F_FD8*2R58IH04E-2_/8OHEFOIC_HE802RR+5mAmph q'#bF5FLFD2_IR5*RI0H8E2-4/OI_EOFHCH_I820ER4+R;F
OMN#0M80RCEb0_lMk_DOCD:#RR0HMCsoCRR:=5mAmph q'#bF5FLFD2_8R8*5CEb0-/428E_OFCHO_b8C0RE2+AR5m mpqbh'FL#5F_FDI*2RRC58b-0E4I2/_FOEH_OC80CbE+2RR
4;0C$bR0Fk_#Lk4$_0bHCR#sRNsRN$5b8C0ME_kOl_C#DD-84RF0IMF,RjR8IH0ME_kOl_C#DD-84RF0IMF2RjRRFV#_08DHFoO#;
HNoMDFRskL0_kR#4:kRF0k_L#04_$;bCRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-.-R7sRNsRN$FsVR_k8F0HR5M0bkRR0F0-sH#00NC
#2#MHoNIDRF_k0L4k#RF:RkL0_k_#40C$b;$
0bFCRkL0_k_#.0C$bRRH#NNss$8R5CEb0_lMk_DOCD4#-RI8FMR0Fj.,R*8IH0ME_kOl_C#DD+84RF0IMF2RjRRFV#_08DHFoO#;
HNoMDFRskL0_kR#.:kRF0k_L#0._$;bCRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-.-R7sRNsRN$FsVR_k8F0HR5M0bkRR0F0-sH#00NC
#2#MHoNIDRF_k0L.k#RF:RkL0_k_#.0C$b;$
0bFCRkL0_k_#c0C$bRRH#NNss$8R5CEb0_lMk_DOCD4#-RI8FMR0Fjc,R*8IH0ME_kOl_C#DD+8dRF0IMF2RjRRFV#_08DHFoO#;
HNoMDFRskL0_kR#c:kRF0k_L#0c_$;bCRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-.-R7sRNsRN$FsVR_k8F0HR5M0bkRR0F0-sH#00NC
#2#MHoNIDRF_k0Lck#RF:RkL0_k_#c0C$b;$
0bFCRkL0_k_#U0C$bRRH#NNss$8R5CEb0_lMk_DOCD4#-RI8FMR0FjU,R*8IH0ME_kOl_C#DD+8(RF0IMF2RjRRFV#_08DHFoO#;
HNoMDFRskL0_kR#U:kRF0k_L#0U_$;bCRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-.-R7sRNsRN$FsVR_k8F0HR5M0bkRR0F0-sH#00NC
#2#MHoNIDRF_k0LUk#RF:RkL0_k_#U0C$b;$
0bbCRN0sH$k_L#0U_$RbCHN#Rs$sNRC58b_0EM_klODCD#R-48MFI0jFR,HRI8_0EM_klODCD#R-48MFI0jFR2VRFR8#0_oDFH
O;#MHoNsDRbHNs0L$_kR#U:NRbs$H0_#LkU$_0bRC;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--.N7Rs$sNRRFVsF_8k50RHkMb0FR0RH0s-N#002C#
o#HMRNDIsbNH_0$LUk#Rb:RN0sH$k_L#0U_$;bC
b0$CkRF0k_L#_4n0C$bRRH#NNss$8R5CEb0_lMk_DOCD4#-RI8FMR0Fj4,RnH*I8_0EM_klODCD#6+4RI8FMR0FjF2RV0R#8F_Do;HO
o#HMRNDs0Fk_#Lk4:nRR0Fk_#Lk40n_$;bCRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-.-R7sRNsRN$FsVR_k8F0HR5M0bkRR0F0-sH#00NC
#2#MHoNIDRF_k0L4k#nRR:F_k0L4k#n$_0b
C;0C$bRsbNH_0$L4k#n$_0bHCR#sRNsRN$5b8C0ME_kOl_C#DD-84RF0IMF,RjRI.*HE80_lMk_DOCD4#+RI8FMR0FjF2RV0R#8F_Do;HO
o#HMRNDssbNH_0$L4k#nRR:bHNs0L$_kn#4_b0$CR;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RR.7NNss$VRFR8s_FRk05bHMk00RFsR0H0-#N#0C2H
#oDMNRNIbs$H0_#Lk4:nRRsbNH_0$L4k#n$_0b
C;0C$bR0Fk_#Lkd0._$RbCHN#Rs$sNRC58b_0EM_klODCD#R-48MFI0jFR,.Rd*8IH0ME_kOl_C#DD+Rd48MFI0jFR2VRFR8#0_oDFH
O;#MHoNsDRF_k0Ldk#.RR:F_k0Ldk#.$_0bRC;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-7R.RsNsNF$RV_Rs80FkRM5HbRk000FRs#H-0CN0##2
HNoMDFRIkL0_k.#dRF:RkL0_k.#d_b0$C0;
$RbCbHNs0L$_k.#d_b0$C#RHRsNsN5$R80CbEk_MlC_OD-D#4FR8IFM0RRj,cH*I8_0EM_klODCD#R+d8MFI0jFR2VRFR8#0_oDFH
O;#MHoNsDRbHNs0L$_k.#dRb:RN0sH$k_L#_d.0C$b;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--.N7Rs$sNRRFVsF_8k50RHkMb0FR0RH0s-N#002C#
o#HMRNDIsbNH_0$Ldk#.RR:bHNs0L$_k.#d_b0$C#;
HNoMDFRskC0_MRR:#_08DHFoOC_POs0F5b8C0ME_kOl_C#DD-84RF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RNCML#DCRsVFRH0s-N#00
C##MHoNIDRF_k0C:MRR8#0_oDFHPO_CFO0sC58b_0EM_klODCD#R-48MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-MRCNCLD#FRVssR0H0-#N#0C
o#HMRNDI_s0C:MRR8#0_oDFHPO_CFO0sC58b_0EM_klODCD#R-48MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-sRIHR0CCLMNDRC#VRFsCENORIsFRRFV)RqvODCD#H
#oDMNR_HMsRCo:0R#8F_Do_HOP0COFIs5HE80+Rd68MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--k8#CRR0FsHCo#s0CRh7QRH
#oDMNRksF0C_soRR:#_08DHFoOC_POs0F58IH0dE+6FR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RCk#8FR0RosCHC#0smR7z#a
HNoMDFRIks0_C:oRR8#0_oDFHPO_CFO0sH5I8+0Ed86RF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-#RkC08RFCRso0H#C7sRm
za#MHoNsDRF_k0s4CoR#:R0D8_FOoH_OPC05FsI0H8ER-48MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-#RkC08RFEROFCF#R0LCIMCCRh7QR8NMR0FkbRk0FAVRD	FORv)q
o#HMRNDs_N8sRCo:0R#8F_Do_HOP0COFNs58I8sHE80-84RF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-k-R#RC80sFRC#oH0RCs)7q7)H
#oDMNR8IN_osCR#:R0D8_FOoH_OPC05FsNs88I0H8ER-48MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--k8#CRR0FsHCo#s0CR7Wq7#)
HNoMDFRDIN_s8R8s:0R#8F_Do_HOP0COF4s5dFR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-NRs8R8sL#H0RbHMk00RFqR)vCRODRD#5LcRHR0#skCJH8sC2H
#oDMNRIDF_8IN8:sRR8#0_oDFHPO_CFO0sd54RI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-R8IN8LsRHR0#HkMb0FR0Rv)qRDOCD5#RcHRL0s#RCHJks2C8
o#HMRND)7q7)l_0bRR:#_08DHFoOC_POs0F58N8s8IH04E-RI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RCk#8FR0RbbHCMDHCqR)7
7)#MHoNWDRq)77_b0lR#:R0D8_FOoH_OPC05FsNs88I0H8ER-48MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--k8#CRR0FbCHbDCHMR7Wq7#)
HNoMDQR7hl_0bRR:#_08DHFoOC_POs0F58IH04E-RI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-k-R#RC80bFRHDbCHRMC7
Qh#MHoNWDR l_0bRR:#_08DHFoOR;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--k8#CRR0FbCHbDCHMR
W #MHoNsDR_8N8sC_soRR:#_08DHFoOC_POs0F58N8s8IH04E-RI8FMR0Fj
2;-C-RML8RD	FORlsNRbHlDCClM00NHRFM#MHoN
D#-L-RCMoHRD#CCRO0sRNlHDlbCMlC0HN0F#MRHNoMDV#
k0MOHRFMo_C0M_kln8c5CEb0:MRH0CCoss2RCs0kMMRH0CCos#RH
sPNHDNLCNRPDRR:HCM0oRCs:j=R;C
Lo
HMRNRPD=R:Rb8C0nE/cR;
RRHV5C58bR0ElRF8nRc2>URc2ER0CRM
RPRRN:DR=NRPDRR+4R;
R8CMR;HV
sRRCs0kMNRPDC;
Mo8RCM0_knl_cV;
k0MOHRFMo_C0D0CVFsPC_5d.80CbERR:HCM0o2CsR0sCkRsMHCM0oRCsHL#
CMoH
sRRCs0kMC58bR0ElRF8n;c2
8CMR0oC_VDC0CFPs._d;k
VMHO0FoMRCD0_CFV0P5Cs80CbERR:HCM0o;CsRGlNRH:RMo0CCRs2skC0sHMRMo0CCHsR#N
PsLHNDPCRN:DRR0HMCsoCRR:=jL;
CMoH
HRRV8R5CEb0Rl-RN>GR=2RjRC0EMR
RRNRPD=R:Rb8C0-ERRGlN;R
RCCD#
RRRRDPNRR:=80CbER;
R8CMR;HV
sRRCs0kMN5PD
2;CRM8o_C0D0CVFsPC;k
VMHO0FoMRCM0_kdl_.C58bR0E:MRH0CCoss2RCs0kMMRH0CCos#RH
sPNHDNLCNRPDRR:HCM0oRCs:j=R;C
Lo
HMRVRHRC58bR0E<c=RUMRN8CR8bR0E>nR42ER0CRM
RRRRPRND:4=R;R
RCRM8H
V;RCRs0MksRDPN;M
C8CRo0k_Ml._d;k
VMHO0FoMRCM0_k4l_nC58bR0E:MRH0CCoss2RCs0kMMRH0CCos#RH
sPNHDNLCNRPDRR:HCM0oRCs:j=R;C
Lo
HMRVRHRC58bR0E<4=RnMRN8CR8bR0E>2RjRC0EMR
RRPRRN:DR=;R4
CRRMH8RVR;
R0sCkRsMP;ND
8CMR0oC_lMk_;4n
MOF#M0N0kRMlC_ODnD_cRR:HCM0oRCs:o=RCM0_knl_cC58b20E;F
OMN#0MD0RCFV0P_Csd:.RR0HMCsoCRR:=o_C0D0CVFsPC_5d.80CbE
2;O#FM00NMRlMk_DOCD._dRH:RMo0CC:sR=CRo0k_Ml._d5VDC0CFPs._d2O;
F0M#NRM0D0CVFsPC_R4n:MRH0CCos=R:R0oC_VDC0CFPsC5DVP0FCds_.d,R.
2;O#FM00NMRlMk_DOCDn_4RH:RMo0CC:sR=CRo0k_Mln_45VDC0CFPsn_42
;
0C$bR0Fk_#Lk_b0$Cc_n##RHRsNsN5$RM_klODCD_Rnc8MFI0jFR,HRI8-0E4FR8IFM0RRj2F#VR0D8_FOoH;$
0bFCRkL0_k0#_$_bCdR.#HN#Rs$sNRk5MlC_ODdD_.FR8IFM0RRj,I0H8ER-48MFI0jFR2VRFR8#0_oDFH
O;0C$bR0Fk_#Lk_b0$Cn_4##RHRsNsN5$RM_klODCD_R4n8MFI0jFR,HRI8-0E4FR8IFM0RRj2F#VR0D8_FOoH;H
#oDMNRksF0k_L#c_n#RR:F_k0L_k#0C$b_#nc;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--.N7Rs$sNRRFV80FkRM5HbRk000FRs#H-0CN0##2
HNoMDFRIkL0_kn#_c:#RR0Fk_#Lk_b0$Cc_n#R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RR.7NNss$VRFRk8F0HR5M0bkRR0F0-sH#00NC
#2#MHoNsDRF_k0L_k#dR.#:kRF0k_L#$_0bdC_.R#;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-7R.RsNsNF$RVFR8k50RHkMb0FR0RH0s-N#002C#
o#HMRNDI0Fk_#Lk_#d.RF:RkL0_k0#_$_bCd;.#
o#HMRNDs0Fk_#Lk_#4nRF:RkL0_k0#_$_bC4;n#RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-.-R7sRNsRN$F8VRFRk05bHMk00RFsR0H0-#N#0C2H
#oDMNRkIF0k_L#n_4#RR:F_k0L_k#0C$b_#4n;H
#oDMNRksF0M_C_:#RR8#0_oDFHPO_CFO0sk5MlC_ODnD_cFR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--CLMNDRC#VRFs0-sH#00NC##
HNoMDFRIkC0_MR_#:0R#8F_Do_HOP0COFMs5kOl_C_DDn8cRF0IMF2Rj;H
#oDMNRksF0M_C_Rd.:0R#8F_Do;HO
o#HMRNDI0Fk__CMd:.RR8#0_oDFH
O;#MHoNsDRF_k0C4M_nRR:#_08DHFoO#;
HNoMDFRIkC0_Mn_4R#:R0D8_FOoH;H
#oDMNR0Is__CM#RR:#_08DHFoOC_POs0F5lMk_DOCDc_nRI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-I-RsCH0RNCML#DCRsVFROCNEFRsIVRFRv)qRDOCD##
HNoMDsRI0M_C_Rd.:0R#8F_Do;HO
o#HMRNDI_s0C4M_nRR:#_08DHFoO#;
HNoMDMRH_osC_:#RR8#0_oDFHPO_CFO0sH5I8-0E4FR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-#RkC08RFCRso0H#C7sRQ
hR#MHoNsDRF_k0s_Co#RR:#_08DHFoOC_POs0F58IH04E-RI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--k8#CRR0FsHCo#s0CRz7maH
#oDMNRkIF0C_soR_#:0R#8F_Do_HOP0COFIs5HE80-84RF0IMF2Rj;RRR
o#HMRNDs_N8s_Co#RR:#_08DHFoOC_POs0F58N8s8IH04E-RI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RCk#8FR0RosCHC#0s7Rq7#)
HNoMDNRI8C_soR_#:0R#8F_Do_HOP0COFNs58I8sHE80-84RF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-k-R#RC80sFRC#oH0RCsq)77
o#HMRNDD_FIs8N8sR_#:0R#8F_Do_HOP0COF6s5RI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-R8N8sHRL0H#RM0bkRR0F)RqvODCD#cR5R0LH#CRsJskHC
82#MHoNDDRFII_Ns88_:#RR8#0_oDFHPO_CFO0sR568MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--Ns88R0LH#MRHbRk00)FRqOvRC#DDRR5cL#H0RJsCkCHs8-2
-MRC8CR#D0CORlsNRbHlDCClM00NHRFM#MHoN
D#Ns00H0LkC3R\s_NlF#VVCR0\:0R#soHM;L

CMoH
zRRcRd:H5VRs8N8sC_soo2RCsMCNR0C-o-RCsMCNR0CLODF	NRslR
RR-R-RRQVNs88I0H8ERR<OHEFOIC_HE80R#N#HRoM'Rj'0kFRMCk#8HRL0R#
RzRRj:RRRRHV58N8s8IH0=ERRR42oCCMsCN0
RSRRFRDIN_s8R8s<"=Rjjjjjjjjjjjjj&"RR8sN_osC5;j2
RSRRFRDIN_I8R8s<"=Rjjjjjjjjjjjjj&"RR8IN_osC5;j2
MSC8CRoMNCs0zCRjR;
RzRR4:RRRRHV58N8s8IH0=ERRR.2oCCMsCN0
DSSFsI_Ns88RR<="jjjjjjjjjjjj&"RR8sN_osC584RF0IMF2Rj;R
SRDRRFII_Ns88RR<="jjjjjjjjjjjj&"RR8IN_osC584RF0IMF2Rj;C
SMo8RCsMCNR0Cz
4;RRRRzR.R:VRHR85N8HsI8R0E=2RdRMoCC0sNCS
SD_FIs8N8s=R<Rj"jjjjjjjjjj&"RR8sN_osC58.RF0IMF2Rj;R
SRDRRFII_Ns88RR<="jjjjjjjjjjj"RR&I_N8s5Co.FR8IFM0R;j2
MSC8CRoMNCs0zCR.R;
RzRRd:RRRRHV58N8s8IH0=ERRRc2oCCMsCN0
DSSFsI_Ns88RR<="jjjjjjjj"jjRs&RNs8_Cdo5RI8FMR0Fj
2;SRRRRIDF_8IN8<sR=jR"jjjjjjjjj&"RR8IN_osC58dRF0IMF2Rj;C
SMo8RCsMCNR0Cz
d;RRRRzRcR:VRHR85N8HsI8R0E=2R6RMoCC0sNCR
SRDRRFsI_Ns88RR<="jjjjjjjjRj"&NRs8C_soR5c8MFI0jFR2S;
RRRRD_FII8N8s=R<Rj"jjjjjj"jjRI&RNs8_Cco5RI8FMR0Fj
2;S8CMRMoCC0sNCcRz;R
RR6RzRRR:H5VRNs88I0H8ERR=no2RCsMCN
0CSRRRRIDF_8sN8<sR=jR"jjjjj"jjRs&RNs8_C6o5RI8FMR0Fj
2;SFSDIN_I8R8s<"=Rjjjjjjjj"RR&I_N8s5Co6FR8IFM0R;j2
MSC8CRoMNCs0zCR6R;
RzRRn:RRRRHV58N8s8IH0=ERRR(2oCCMsCN0
RSRRFRDIN_s8R8s<"=Rjjjjj"jjRs&RNs8_Cno5RI8FMR0Fj
2;SFSDIN_I8R8s<"=Rjjjjj"jjRI&RNs8_Cno5RI8FMR0Fj
2;S8CMRMoCC0sNCnRz;R
RR(RzRRR:H5VRNs88I0H8ERR=Uo2RCsMCN
0CSRRRRIDF_8sN8<sR=jR"jjjjj&"RR8sN_osC58(RF0IMF2Rj;S
SD_FII8N8s=R<Rj"jjjjj"RR&I_N8s5Co(FR8IFM0R;j2
MSC8CRoMNCs0zCR(R;
RzRRU:RRRRHV58N8s8IH0=ERRRg2oCCMsCN0
RSRRFRDIN_s8R8s<"=Rjjjjj&"RR8sN_osC58URF0IMF2Rj;S
SD_FII8N8s=R<Rj"jj"jjRI&RNs8_CUo5RI8FMR0Fj
2;S8CMRMoCC0sNCURz;R
RRgRzRRR:H5VRNs88I0H8ERR=4Rj2oCCMsCN0
RSRRFRDIN_s8R8s<"=Rjjjj"RR&s_N8s5CogFR8IFM0R;j2
DSSFII_Ns88RR<="jjjj&"RR8IN_osC58gRF0IMF2Rj;C
SMo8RCsMCNR0Cz
g;RRRRzR4jRH:RVNR58I8sHE80R4=R4o2RCsMCN
0CSRRRRIDF_8sN8<sR=jR"jRj"&NRs8C_soj54RI8FMR0Fj
2;SFSDIN_I8R8s<"=Rj"jjRI&RNs8_C4o5jFR8IFM0R;j2
MSC8CRoMNCs0zCR4
j;RRRRzR44RH:RVNR58I8sHE80R4=R.o2RCsMCN
0CSRRRRIDF_8sN8<sR=jR"j&"RR8sN_osC5R448MFI0jFR2S;
SIDF_8IN8<sR=jR"j&"RR8IN_osC5R448MFI0jFR2S;
CRM8oCCMsCN0R4z4;R
RR4Rz.:RRRRHV58N8s8IH0=ERR24dRMoCC0sNCR
SRDRRFsI_Ns88RR<='Rj'&NRs8C_so.54RI8FMR0Fj
2;SFSDIN_I8R8s<'=Rj&'RR8IN_osC5R4.8MFI0jFR2S;
CRM8oCCMsCN0R.z4;R
RR4Rzd:RRRRHV58N8s8IH0>ERR24dRMoCC0sNCR
SRDRRFsI_Ns88RR<=s_N8s5Co48dRF0IMF2Rj;R
SRDRRFII_Ns88RR<=I_N8s5Co48dRF0IMF2Rj;C
SMo8RCsMCNR0Cz;4d
R
RR-R-RRQV5M8H_osC2CRso0H#C7sRQkhR#oHMRiBp
RRRRcz4RRR:H5VR8_HMs2CoRMoCC0sNCR
RRRRRRsRbF#OC#BR5pRi,72QhRoLCHRM
RRRRRRRRRHRRVBR5p=iRR''4R8NMRiBp'CCPMR020MEC
RRRRRRRRRRRRRRRR_HMsRCo<5=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj&"RRh7Q2R;
RRRRRRRRRCRRMH8RVR;
RRRRRCRRMb8RsCFO#
#;S8CMRMoCC0sNC4RzcR;
RzRR4R6R:VRHRF5M0HR8MC_soo2RCsMCN
0CRRRRRRRRRRRRHsM_C<oR="R5jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"RR&72Qh;C
SMo8RCsMCNR0Cz;46
R
RR-R-RRQV5Fs8ks0_CRo2sHCo#s0CR7)_mRzakM#Ho_R)miBp
RRRRnz4sk8F0:RRRRHV5Fs8ks0_CRo2oCCMsCN0
RRRRRRRRFbsO#C#R_5)miBp,FRsks0_C2o4RoLCHRM
RRRRRRRRRHRRV)R5_pmBiRR='R4'NRM8)B_mpCi'P0CM2ER0CRM
RRRRRRRRRRRRR)RR_z7ma=R<RksF0C_so
4;RRRRRRRRRRRRCRM8H
V;RRRRRRRRCRM8bOsFC;##
RRRRRRRR8CMRMoCC0sNC4RznFs8k
0;RRRRzs4(80FkRRR:H5VRMRF0sk8F0C_soo2RCsMCN
0CRRRRRRRRRRRR)m_7z<aR=FRsks0_C;o4
MSC8CRoMNCs0zCR48(sF;k0
z
S48nIFRk0RH:RVIR580Fk_osC2CRoMNCs0RC
RRRRRbRRsCFO#5#RWB_mpRi,I0Fk_osC2CRLo
HMRRRRRRRRRRRRH5VRWB_mp=iRR''4R8NMRmW_B'piCMPC002RE
CMRRRRRRRRRRRRRRRRWm_7z<aR=FRIks0_CIo5HE80-84RF0IMF2Rj;R
RRRRRRRRRRMRC8VRH;R
RRRRRRMRC8sRbF#OC#R;
RRRRRCRRMo8RCsMCNR0CzI4n80Fk;R
RR4Rz(FI8kR0R:VRHRF5M08RIF_k0s2CoRMoCC0sNCR
RRRRRRRRRR_RW7amzRR<=I0Fk_osC58IH04E-RI8FMR0Fj
2;S8CMRMoCC0sNC4Rz(FI8k
0;
RRRRR--Q5VRs8N8sC_sos2RC#oH0RCs)7q7)#RkHRMomiBp
RRRRnz4s:RRRRHV58sN8ss_CRo2oCCMsCN0
R--RRRRRbRRsCFO#5#RmiBp,qR)727)RoLCH-M
-RRRRRRRRRRRRRHV5pmBiRR='R4'NRM8miBp'CCPMR020MEC
R--RRRRRRRRRRRRRsRRNs8_C<oR=qR)757)Ns88I0H8ER-48MFI0jFR2-;
-RRRRRRRRRRRR8CMR;HV
R--RRRRRCRRMb8RsCFO#
#;-C-SMo8RCsMCNR0Czs4n;-
-RRRRzs4(RH:RVMR5Fs0RNs88_osC2CRoMNCs0RC
RRRRRRRRRsRRNs8_C<oR=qR)7;7)
MSC8CRoMNCs0zCR4;ns
-
S-VRQRN5I8_8ss2CoRosCHC#0sqRW7R7)kM#Ho_RWmiBp
RRRRnz4I:RRRRHV58IN8ss_CRo2oCCMsCN0
RRRRRRRRFbsO#C#Rp5BiW,Rq)772CRLo
HMRRRRRRRRRRRRH5VRBRpi=4R''MRN8pRBiP'CC2M0RC0EMR
RRRRRRRRRRRRRRNRI8C_so=R<R7Wq7N)58I8sHE80-84RF0IMF2Rj;R
RRRRRRRRRRMRC8VRH;R
RRRRRRMRC8sRbF#OC#S;
CRM8oCCMsCN0Rnz4IR;
RzRR4R(I:VRHRF5M0NRI8_8ss2CoRMoCC0sNCR
RRRRRRRRRRNRI8C_so=R<R7Wq7
);S8CMRMoCC0sNC4Rz(
I;
RRRRR-- sG0NFRDoRHOVRFs7DkNRsbF0NRO#SC
-F-M0CRMC88CRsVFR_MFsOI_E	CO
-S-zosCRb:RsCFO#B#5pRi2LHCoM-
-SHRRVBR5p i'ea hR8NMRiBpR'=R4R'20MEC
S--R7RRQ0h_l<bR=QR7h-;
-RSRR7)q70)_l<bR=qR)7;7)
S--RWRRq)77_b0lRR<=W7q7)-;
-RSRR_W 0Rlb<W=R -;
-RSRCRM8H
V;-C-SMb8RsCFO#
#;
-S-RRQV)8CNR8q8s#C#RW=RsCH0R8q8s#C#,$RLb#N#Rh7QRR0FFbk0kH0RV RWRRH#CLMND
C8SkzlGRR:bOsFC5##W0 _lRb,)7q7)l_0bW,Rq)77_b0l,QR7hl_0bs,RF_k0s2Co
RSRLHCoM-
-SRRRRRHV57Wq70)_l=bRR7)q70)_lNbRMW8R l_0bRR='24'RC0EM-
-SRSRs0Fk_osC4=R<Rh7Q_b0l;-
-SDSC#SC
SsRRF_k0s4CoRR<=s0Fk_osC58IH04E-RI8FMR0Fj
2;-S-SCRM8H
V;S8CMRFbsO#C#;R
SR
RRRRRR-t-RCsMCNR0C0REC)RqvODCD#MRN8CR#D0CORoDFHVORF)sRq4vAn4_1_
14SUz4RH:RVOR5EOFHCH_I8R0E=2R4RMoCC0sNCR
SRRSRREzO	H:RVNR58I8sHE80R4>Rco2RCsMCN
0CRRRRRRRRk	ODRb:RsCFO#B#5p
i2RRRRRRRRRoLCHRM
RRRRRRRRRRHV5iBp'CCPMN0RMB8Rp=iRR''42ER0CRM
RRRRRRRRRsRR_8N8sC_so85N8HsI8-0E4FR8IFM0R24cRR<=)7q7)85N8HsI8-0E4FR8IFM0R24c;R
RRRRRRRRRCRM8H
V;RRRRRRRRCRM8bOsFCR##k	OD;R
SR8CMRMoCC0sNCORzE
	;RRRRSgz4RV:RFHsRRRHM5b8C0ME_kOl_C#DDR4-R2FR8IFM0RojRCsMCN
0CSR--Q5VRNs88I0H8ERR>4Rc2M8CCRR0FONsC0ICRsCH0RNCMLRDCNRM8Fbk0kC0RMDNLCCR#D0CORoDFHRO
RRRRRSRRzR.j:VRHR85N8HsI8R0E>cR42CRoMNCs0SC
-V-RHVGRFOsRNRDD4UdU(#,RCODC0VRFRH0s#00NCFRM0CRLHRMosHCo#s0CCS8
SsSSF_k0CHM52=R<R''4RCIEMsR5_8N8sC_so85N8HsI8-0E4FR8IFM0R24cRH=R2DRC#'CRj
';SSSSI0Fk_5CMH<2R=4R''ERIC5MRI_N8s5CoNs88I0H8ER-48MFI04FRc=2RRRH2CCD#R''j;R
RRRRRRRRRRRRRRsRI0M_C5RH2<W=R ERIC5MRI_N8s5CoNs88I0H8ER-48MFI04FRc=2RRRH2CCD#R''j;R
RRRRRRCRSMo8RCsMCNR0Cz;.j
-S-RRQV58N8s8IH0<ER=cR42FRMRHIs0CCRMDNLCsRFR0FkbRk0CLMND#CRCODC0FRDoRHOM8CCCR8
SRRRR.Sz4RR:H5VRNs88I0H8E=R<R24cRMoCC0sNCS
SSFSskC0_M25HRR<=';4'
SSSSkIF0M_C5RH2<'=R4
';RRRRRRRRRRRRRRRRI_s0CHM52=R<R;W 
RRRRRRRRMSC8CRoMNCs0zCR.
4;SR--tCCMsCN0RC0ERv)qRDOCDN#RM08Rs#H-0CN0#R
RRRRRRzRS.:.RRsVFRH[RMIR5HE80_lMk_DOCD-#RRR428MFI0jFRRMoCC0sNCR
RRRRRRRRRRRRRR0RN0LsHkR0C\N3slV_FV0#C\VRFRqA)vn_4dXUc4:7RRLDNCHDR#WR""R;
RRRRRRRRRRRRRLRRCMoH
RRRRRRRRRRRR)SAq4v_ncdUXR47:qR)vnA4__141S4
RRRRRRRRRRRRb0FsRblNRQ57q25jRR=>HsM_C[o52q,R7q7)RR=>D_FII8N8sd54RI8FMR0FjR2,7RQA=">RjR",q)77A>R=RIDF_8sN84s5dFR8IFM0R,j2
SSSSq hRR=>',4'R)11q>R=R''j, RWq>R=R0Is_5CMHR2,BqpiRR=>B,piRA hRR=>',4'R)11A>R=R''j, RWA>R=R''j,pRBi=AR>pRBiS,
SRSRRmR7q25jRR=>I0Fk_#Lk4,5H[R2,75mAj=2R>FRskL0_k5#4H2,[2
;
RRRRRRRRRRRRRRRRs0Fk_osC5R[2<s=RF_k0L4k#5[H,2ERIC5MRs0Fk_5CMH=2RR''42DRC#'CRZ
';SSSSI0Fk_osC5R[2<I=RF_k0L4k#5KH,2ERIC5MRI0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRS8CMRMoCC0sNC.Rz.R;
RRRRS8CMRMoCC0sNC4RzgR;
RCRRMo8RCsMCNR0Cz;4URRRR
RRRR
RRRRRR-t-RCsMCNR0C0REC)RqvODCD#MRN8CR#D0CORoDFHVORF)sRq4vAn._1_
1.Sdz.RH:RVOR5EOFHCH_I8R0E=2R.RMoCC0sNCR
SREzO	RR:H5VRNs88I0H8ERR>4Rd2oCCMsCN0
RRRRRRRRDkO	RR:bOsFC5##B2pi
RRRRRRRRCRLo
HMRRRRRRRRRVRHRp5BiP'CCRM0NRM8BRpi=4R''02RE
CMRRRRRRRRRRRRs8_N8ss_CNo58I8sHE80-84RF0IMFdR42=R<R7)q7N)58I8sHE80-84RF0IMFdR42R;
RRRRRRRRR8CMR;HV
RRRRRRRR8CMRFbsO#C#RDkO	S;
RMRC8CRoMNCs0zCRO;E	
RRRR.SzcRR:VRFsHMRHRC58b_0EM_klODCD#RR-482RF0IMFRRjoCCMsCN0
-S-RRQV58N8s8IH0>ERR24dRCMC8FR0RCOsNR0CI0sHCMRCNCLDR8NMR0FkbRk0CLMND#CRCODC0FRDo
HORRRRRRRRS6z.RH:RVNR58I8sHE80R4>Rdo2RCsMCN
0CSR--VRHGVRFsODNDRU4dUR(,#CCDOF0RVsR0HN#00MCRFL0RCoHMRosCHC#0s
C8RRRRRRRRRRRRRRRRs0Fk_5CMH<2R=4R''ERIC5MRs8_N8ss_CNo58I8sHE80-84RF0IMFdR42RR=HC2RDR#C';j'
SSSSkIF0M_C5RH2<'=R4I'RERCM58IN_osC58N8s8IH04E-RI8FMR0F4Rd2=2RHR#CDCjR''R;
RRRRRRRRRRRRRIRRsC0_M25HRR<=WI RERCM58IN_osC58N8s8IH04E-RI8FMR0F4Rd2=2RHR#CDCjR''R;
RRRRRSRRCRM8oCCMsCN0R6z.;-
S-VRQR85N8HsI8R0E<4=RdM2RFsRIHR0CCLMNDFCRskRF00bkRNCMLRDC#CCDOD0RFOoHRCMC8
C8RRSRRzRS.:nRRRHV58N8s8IH0<ER=dR42CRoMNCs0SC
RRRRRRRRRRRRs0Fk_5CMH<2R=4R''S;
SISSF_k0CHM52=R<R''4;R
RRRRRRRRRRRRRRsRI0M_C5RH2<W=R R;
RRRRRSRRCRM8oCCMsCN0Rnz.;-
S-CRtMNCs00CRE)CRqOvRC#DDR8NMRH0s-N#00
C#RRRRRRRRS(z.RV:RF[sRRRHM58IH0ME_kOl_C#DDR4-R2FR8IFM0RojRCsMCN
0CRRRRRRRRRRRRRRRRNs00H0LkC3R\s_NlF#VVCR0\FAVR)_qvU.4gXR.7:NRDLRCDH"#RW
";RRRRRRRRRRRRRRRRLHCoMR
RRRRRRRRRRARS)_qvU.4gXR.7:qR)vnA4__1.1S.
RRRRRRRRRRRRb0FsRblNRQ57q>R=R_HMs5Co.+*[4FR8IFM0R[.*2q,R7q7)RR=>D_FII8N8s.54RI8FMR0FjR2,7RQA=">Rj,j"R7q7)=AR>FRDIN_s858s48.RF0IMF2Rj,S
SSRRRRq hRR=>',4'R)11q>R=R''j, RWq>R=R0Is_5CMHR2,BqpiRR=>B,piRA hRR=>',4'R)11A>R=R''j, RWA>R=R''j,pRBi=AR>pRBiS,
SRSRRmR7q254RR=>I0Fk_#Lk.,5H.+*[4R2,75mqj=2R>FRIkL0_k5#.H*,.[R2,75mA4=2R>FRskL0_k5#.H*,.[2+4,mR7A25jRR=>s0Fk_#Lk.,5HR[.*2
2;RRRRRRRRRRRRRRRRs0Fk_osC5[.*2=R<RksF0k_L#H.5,[.*2ERIC5MRs0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRs0Fk_osC5[.*+R42<s=RF_k0L.k#5.H,*4[+2ERIC5MRs0Fk_5CMH=2RR''42DRC#'CRZ
';SSSSI0Fk_osC5[.*2=R<RkIF0k_L#H.5,[.*2ERIC5MRI0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRI0Fk_osC5[.*+R42<I=RF_k0L.k#5.H,*4[+2ERIC5MRI0Fk_5CMH=2RR''42DRC#'CRZ
';
RRRRRRRRMSC8CRoMNCs0zCR.
(;RRRRRMSC8CRoMNCs0zCR.
c;RRRRCRM8oCCMsCN0Rdz.;
RR
RSRR-R-RMtCC0sNCER0CqR)vCRODRD#NRM8#CCDOD0RFOoHRsVFRv)qA_4n11c_cz
S.:URRRHV5FOEH_OCI0H8ERR=co2RCsMCN
0CSEzO	H:RVNR58I8sHE80R4>R.o2RCsMCNR0C
RRRRRRRRDkO	RR:bOsFC5##B2pi
RRRRRRRRCRLo
HMRRRRRRRRRVRHRp5BiP'CCRM0NRM8BRpi=4R''02RE
CMRRRRRRRRRRRRs8_N8ss_CNo58I8sHE80-84RF0IMF.R42=R<R7)q7N)58I8sHE80-84RF0IMF.R42R;
RRRRRRRRR8CMR;HV
RRRRRRRR8CMRFbsO#C#RDkO	S;
RMRC8CRoMNCs0zCRO;E	
RRRR.SzgRR:VRFsHMRHRC58b_0EM_klODCD#RR-482RF0IMFRRjoCCMsCN0
-S-RRQV58N8s8IH0>ERR24.RCMC8FR0RCOsNR0CI0sHCMRCNCLDR8NMR0FkbRk0CLMND#CRCODC0FRDo
HORRRRRRRRSjzdRH:RVNR58I8sHE80R4>R.o2RCsMCN
0CSR--VRHGVRFsODNDRU4dUR(,#CCDOF0RVsR0HN#00MCRFL0RCoHMRosCHC#0s
C8RRRRRRRRRRRRRRRRs0Fk_5CMH<2R=4R''ERIC5MRs8_N8ss_CNo58I8sHE80-84RF0IMF.R42RR=HC2RDR#C';j'
SSSSkIF0M_C5RH2<'=R4I'RERCM58IN_osC58N8s8IH04E-RI8FMR0F4R.2-2RHR#CDCjR''R;
RRRRRRRRRRRRRIRRsC0_M25HRR<=WI RERCM58IN_osC58N8s8IH04E-RI8FMR0F4R.2=2RHR#CDCjR''R;
RRRRRSRRCRM8oCCMsCN0Rjzd;-
S-VRQR85N8HsI8R0E<4=R.M2RFsRIHR0CCLMNDFCRskRF00bkRNCMLRDC#CCDOD0RFOoHRCMC8
C8RRSRRzRSd:4RRRHV58N8s8IH0<ER=.R42CRoMNCs0SC
SsSSF_k0CHM52=R<R''4;S
SSFSIkC0_M25HRR<=';4'
RRRRRRRRRRRRRRRR0Is_5CMH<2R= RW;R
RRRRRRCRSMo8RCsMCNR0Cz;d4
-S-RMtCC0sNCER0CqR)vCRODRD#NRM80-sH#00NCR#
RRRRRSRRzRd.:FRVsRR[H5MRI0H8Ek_MlC_ODRD#-2R4RI8FMR0FjCRoMNCs0RC
RRRRRRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)RAqcv_jXgnc:7RRLDNCHDR#WR""R;
RRRRRRRRRRRRRLRRCMoH
RRRRRRRRRRRR)SAqcv_jXgnc:7RRv)qA_4n11c_cR
SRRRRRRRRRbRRFRs0lRNb5q7QRR=>HsM_Cco5*d[+RI8FMR0Fc2*[,7Rq7R)q=D>RFII_Ns885R448MFI0jFR27,RQ=AR>jR"j"jj,7Rq7R)A=D>RFsI_Ns885R448MFI0jFR2S,
S SSh=qR>4R''1,R1R)q='>RjR',WR q=I>RsC0_M25H,pRBi=qR>pRBi ,Rh=AR>4R''1,R1R)A='>RjR',WR A='>RjR',BApiRR=>B,pi
SSSSq7m5Rd2=I>RF_k0Lck#5RH,c+*[dR2,
SSSSq7m5R.2=I>RF_k0Lck#5cH,*.[+2
,RSSSS75mq4=2R>FRIkL0_k5#cH*,c[2+4,SR
S7SSmjq52>R=RkIF0k_L#Hc5,*Rc[
2,SSSS75mAd=2R>FRskL0_k5#cHc,R*d[+2
,RSSSS75mA.=2R>FRskL0_k5#cH*,c[2+.,SR
S7SSm4A52>R=RksF0k_L#Hc5,[c*+,42RS
SSmS7A25jRR=>s0Fk_#Lkc,5HR[c*2
2;SSSSs0Fk_osC5[c*2=R<RksF0k_L#Hc5,[c*2ERIC5MRs0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRs0Fk_osC5[c*+R42<s=RF_k0Lck#5cH,*4[+2ERIC5MRs0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRs0Fk_osC5[c*+R.2<s=RF_k0Lck#5cH,*.[+2ERIC5MRs0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRs0Fk_osC5[c*+Rd2<s=RF_k0Lck#5cH,*d[+2ERIC5MRs0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRI0Fk_osC5[c*2=R<RkIF0k_L#Hc5,[c*2ERIC5MRI0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRI0Fk_osC5[c*+R42<I=RF_k0Lck#5cH,*4[+2ERIC5MRI0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRI0Fk_osC5[c*+R.2<I=RF_k0Lck#5cH,*.[+2ERIC5MRI0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRI0Fk_osC5[c*+Rd2<I=RF_k0Lck#5cH,*d[+2ERIC5MRI0Fk_5CMH=2RR''42DRC#'CRZ
';
RRRRRRRRMSC8CRoMNCs0zCRd
.;RRRRRMSC8CRoMNCs0zCR.
g;RRRRCRM8oCCMsCN0RUz.;S

RRRR-t-RCsMCNR0C0REC)RqvODCD#MRN8CR#D0CORoDFHVORF)sRq4vAng_1_
1gSdzdRH:RVOR5EOFHCH_I8R0E=2RgRMoCC0sNCz
SORE	:VRHR85N8HsI8R0E>4R42CRoMNCs0RC
RRRRRkRRORD	:sRbF#OC#p5BiR2
RRRRRRRRLHCoMR
RRRRRRRRRH5VRB'piCMPC0MRN8pRBiRR='24'RC0EMR
RRRRRRRRRR_RsNs88_osC58N8s8IH04E-RI8FMR0F4R42<)=Rq)7758N8s8IH04E-RI8FMR0F4;42
RRRRRRRRCRRMH8RVR;
RRRRRCRRMb8RsCFO#k#RO;D	
RSRCRM8oCCMsCN0REzO	R;
RSRRzRdc:FRVsRRHH5MR80CbEk_MlC_ODRD#-2R4RI8FMR0FjCRoMNCs0SC
-Q-RVNR58I8sHE80R4>R4M2RCRC80OFRs0CNCsRIHR0CCLMNDNCRMF8Rkk0b0MRCNCLDRD#CCRO0DHFoOR
RRRRRRzRSd:6RRRHV58N8s8IH0>ERR244RMoCC0sNC-
S-HRVGFRVsNROD4DRd(UU,CR#D0CORRFV0#sH0CN0R0MFRHLCMsoRC#oH0CCs8R
RRRRRRRRRRRRRRFRskC0_M25HRR<='R4'IMECR_5sNs88_osC58N8s8IH04E-RI8FMR0F4R42=2RHR#CDCjR''S;
SISSF_k0CHM52=R<R''4RCIEMIR5Ns8_CNo58I8sHE80-84RF0IMF4R42RR=HC2RDR#C';j'
RRRRRRRRRRRRRRRR0Is_5CMH<2R= RWRCIEMIR5Ns8_CNo58I8sHE80-84RF0IMF4R42RR=HC2RDR#C';j'
RRRRRRRRMSC8CRoMNCs0zCRd
6;SR--Q5VRNs88I0H8E=R<R244RRMFI0sHCMRCNCLDRRFsFbk0kC0RMDNLCCR#D0CORoDFHMORCCC88S
RRRRRSnzdRH:RVNR58I8sHE80RR<=4R42oCCMsCN0
RSRRRRRRRRRRFRskC0_M25HRR<=';4'
SSSSkIF0M_C5RH2<'=R4
';RRRRRRRRRRRRRRRRI_s0CHM52=R<R;W 
RRRRRRRRMSC8CRoMNCs0zCRd
n;SR--tCCMsCN0RC0ERv)qRDOCDN#RM08Rs#H-0CN0#R
RRRRRRzRSd:(RRsVFRH[RMIR5HE80_lMk_DOCD-#RRR428MFI0jFRRMoCC0sNCR
RRRRRRRRRRRRRR0RN0LsHkR0C\N3slV_FV0#C\VRFRqA)vj_.cUUX7RR:DCNLD#RHR""W;R
RRRRRRRRRRRRRRCRLo
HMRRRRRRRRRRRRSqA)vj_.cUUX7RR:)Aqv41n_gg_1
RRRRRRRRRRRRRRRRbRRFRs0lRNb5q7QRR=>HsM_Cgo5*([+RI8FMR0Fg2*[,7Rq7R)q=D>RFII_Ns885R4j8MFI0jFR27,RQ=AR>jR"jjjjj"jj,7Rq7R)A=D>RFsI_Ns885R4j8MFI0jFR2S,
S SSh=qR>4R''1,R1R)q='>RjR',WR q=I>RsC0_M25H,pRBi=qR>pRBi ,Rh=AR>4R''1,R1R)A='>RjR',WR A='>RjR',BApiRR=>B,piRS
SSmS7q25(RR=>I0Fk_#LkU,5HU+*[(R2,
SSSSq7m5Rn2=I>RF_k0LUk#5UH,*n[+2
,RSSSS75mq6=2R>FRIkL0_k5#UH*,U[2+6,SR
S7SSmcq52>R=RkIF0k_L#HU5,[U*+,c2RS
SSmS7q25dRR=>I0Fk_#LkU,5HU+*[dR2,
SSSSq7m5R.2=I>RF_k0LUk#5UH,*.[+2
,RSSSS75mq4=2R>FRIkL0_k5#UH*,U[2+4,SR
S7SSmjq52>R=RkIF0k_L#HU5,[U*2
,RSSSS75mA(=2R>FRskL0_k5#UH*,U[2+(,SR
S7SSmnA52>R=RksF0k_L#HU5,[U*+,n2RS
SSmS7A256RR=>s0Fk_#LkU,5HU+*[6R2,
SSSSA7m5Rc2=s>RF_k0LUk#5UH,*c[+2
,RSSSS75mAd=2R>FRskL0_k5#UH*,U[2+d,SR
S7SSm.A52>R=RksF0k_L#HU5,[U*+,.2RS
SSmS7A254RR=>s0Fk_#LkU,5HU+*[4R2,
SSSSA7m5Rj2=s>RF_k0LUk#5UH,*,[2RR
RRRRRRRRRRRRRRRRRRRRRRRRRRQR7ujq52>R=R_HMs5Cog+*[UR2,7AQuRR=>",j"
RRRRRRRRRRRRRRRRRRRRRRRRRRRRu7mq25jRR=>IsbNH_0$LUk#5[H,27,Rm5uAj=2R>bRsN0sH$k_L#HU5,2[2;R
RRRRRRRRRRRRRRFRsks0_Cgo5*R[2<s=RF_k0LUk#5UH,*R[2IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRFRsks0_Cgo5*4[+2=R<RksF0k_L#HU5,[U*+R42IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRFRsks0_Cgo5*.[+2=R<RksF0k_L#HU5,[U*+R.2IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRFRsks0_Cgo5*d[+2=R<RksF0k_L#HU5,[U*+Rd2IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRFRsks0_Cgo5*c[+2=R<RksF0k_L#HU5,[U*+Rc2IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRFRsks0_Cgo5*6[+2=R<RksF0k_L#HU5,[U*+R62IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRFRsks0_Cgo5*n[+2=R<RksF0k_L#HU5,[U*+Rn2IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRFRsks0_Cgo5*([+2=R<RksF0k_L#HU5,[U*+R(2IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRFRsks0_Cgo5*U[+2=R<RNsbs$H0_#LkU,5H[I2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRkIF0C_so*5g[<2R=FRIkL0_k5#UH*,U[I2RERCM5kIF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRkIF0C_so*5g[2+4RR<=I0Fk_#LkU,5HU+*[4I2RERCM5kIF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRkIF0C_so*5g[2+.RR<=I0Fk_#LkU,5HU+*[.I2RERCM5kIF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRkIF0C_so*5g[2+dRR<=I0Fk_#LkU,5HU+*[dI2RERCM5kIF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRkIF0C_so*5g[2+cRR<=I0Fk_#LkU,5HU+*[cI2RERCM5kIF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRkIF0C_so*5g[2+6RR<=I0Fk_#LkU,5HU+*[6I2RERCM5kIF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRkIF0C_so*5g[2+nRR<=I0Fk_#LkU,5HU+*[nI2RERCM5kIF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRkIF0C_so*5g[2+(RR<=I0Fk_#LkU,5HU+*[(I2RERCM5kIF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRkIF0C_so*5g[2+URR<=IsbNH_0$LUk#5[H,2ERIC5MRI0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRS8CMRMoCC0sNCdRz(R;
RRRRS8CMRMoCC0sNCdRzcR;
RCRRMo8RCsMCNR0Cz;dd
R
SR-RR-CRtMNCs00CRE)CRqOvRC#DDR8NMRD#CCRO0DHFoOFRVsqR)vnA4_U14_U14
dSzURR:H5VROHEFOIC_HE80R4=RUo2RCsMCN
0CSEzO	RR:H5VRNs88I0H8ERR>4Rj2oCCMsCN0
RRRRRRRRDkO	RR:bOsFC5##B2pi
RRRRRRRRCRLo
HMRRRRRRRRRVRHRp5BiP'CCRM0NRM8BRpi=4R''02RE
CMRRRRRRRRRRRRs8_N8ss_CNo58I8sHE80-84RF0IMFjR42=R<R7)q7N)58I8sHE80-84RF0IMFjR42R;
RRRRRRRRR8CMR;HV
RRRRRRRR8CMRFbsO#C#RDkO	S;
RCRRMo8RCsMCNR0Cz	OE;R
RRzRSd:gRRsVFRHHRM8R5CEb0_lMk_DOCD-#RRR428MFI0jFRRMoCC0sNC-
S-VRQR85N8HsI8R0E>jR42CRMC08RFsROCCN0RHIs0CCRMDNLCMRN8kRF00bkRNCMLRDC#CCDOD0RFOoH
RRRRRRRRcSzjRR:H5VRNs88I0H8ERR>4Rj2oCCMsCN0
-S-RGVHRsVFRDONDdR4U,U(RD#CCRO0F0VRs0H#NR0CMRF0LMCHoCRso0H#C8sC
RRRRRRRRRRRRRRRRksF0M_C5RH2<'=R4I'RERCM5Ns_8_8ss5CoNs88I0H8ER-48MFI04FRj=2RRRH2CCD#R''j;S
SSFSIkC0_M25HRR<='R4'IMECRN5I8C_so85N8HsI8-0E4FR8IFM0R24jRH=RRC2RDR#C';j'
RRRRRRRRRRRRRRRR0Is_5CMH<2R= RWRCIEMIR5Ns8_CNo58I8sHE80-84RF0IMFjR42RR=HC2RDR#C';j'
RRRRRRRRMSC8CRoMNCs0zCRc
j;SR--Q5VRNs88I0H8E=R<R24jRRMFI0sHCMRCNCLDRRFsFbk0kC0RMDNLCCR#D0CORoDFHMORCCC88S
RRRRRS4zcRH:RVNR58I8sHE80RR<=4Rj2oCCMsCN0
RSRRRRRRRRRRFRskC0_M25HRR<=';4'
SSSSkIF0M_C5RH2<'=R4
';RRRRRRRRRRRRRRRRI_s0CHM52=R<R;W 
RRRRRRRRMSC8CRoMNCs0zCRc
4;SR--tCCMsCN0RC0ERv)qRDOCDN#RM08Rs#H-0CN0#R
RRRRRRzRSc:.RRsVFRH[RMIR5HE80_lMk_DOCD-#RRR428MFI0jFRRMoCC0sNCR
RRRRRRRRRRRRRR0RN0LsHkR0C\N3slV_FV0#C\VRFRqA)vj_4.4cXn:7RRLDNCHDR#WR""R;
RRRRRRRRRRRRRLRRCMoH
RRRRRRRRRRRR)SAq4v_jX.c4Rn7:qR)vnA4_U14_U14
RRRRRRRRRRRRRRRRbRRFRs0lRNb5q7QRR=>HsM_C4o5U+*[486RF0IMFUR4*,[2R7q7)=qR>FRDIN_I858sgFR8IFM0R,j2RA7QRR=>"jjjjjjjjjjjjjjjjR",q)77A>R=RIDF_8sN8gs5RI8FMR0Fj
2,SSSS Rhq='>R4R',1q1)RR=>',j'RqW RR=>I_s0CHM52B,RpRiq=B>RpRi, RhA='>R4R',1A1)RR=>',j'RAW RR=>',j'RiBpA>R=RiBp,SR
S7SSm4q56=2R>FRIkL0_kn#454H,n+*[4,62RS
SSmS7qc542>R=RkIF0k_L#54nHn,4*4[+cR2,
SSSSq7m524dRR=>I0Fk_#Lk4Hn5,*4n[d+42
,RSSSS75mq4R.2=I>RF_k0L4k#n,5H4[n*+24.,SR
S7SSm4q54=2R>FRIkL0_kn#454H,n+*[4,42RS
SSmS7qj542>R=RkIF0k_L#54nHn,4*4[+jR2,
SSSSq7m5Rg2=I>RF_k0L4k#n,5H4[n*+,g2RS
SSmS7q25URR=>I0Fk_#Lk4Hn5,*4n[2+U,SR
S7SSm(q52>R=RkIF0k_L#54nHn,4*([+2
,RSSSS75mqn=2R>FRIkL0_kn#454H,n+*[nR2,
SSSSq7m5R62=I>RF_k0L4k#n,5H4[n*+,62RS
SSmS7q25cRR=>I0Fk_#Lk4Hn5,*4n[2+c,SR
S7SSmdq52>R=RkIF0k_L#54nHn,4*d[+2
,RSSSS75mq.=2R>FRIkL0_kn#454H,n+*[.R2,
SSSSq7m5R42=I>RF_k0L4k#n,5H4[n*+,42RS
SSmS7q25jRR=>I0Fk_#Lk4Hn5,*4n[R2,
SSSSA7m5246RR=>s0Fk_#Lk4Hn5,*4n[6+42
,RSSSS75mA4Rc2=s>RF_k0L4k#n,5H4[n*+24c,SR
S7SSm4A5d=2R>FRskL0_kn#454H,n+*[4,d2RS
SSmS7A.542>R=RksF0k_L#54nHn,4*4[+.R2,
SSSSA7m5244RR=>s0Fk_#Lk4Hn5,*4n[4+42
,RSSSS75mA4Rj2=s>RF_k0L4k#n,5H4[n*+24j,SR
S7SSmgA52>R=RksF0k_L#54nHn,4*g[+2
,RSSSS75mAU=2R>FRskL0_kn#454H,n+*[UR2,
SSSSA7m5R(2=s>RF_k0L4k#n,5H4[n*+,(2RS
SSmS7A25nRR=>s0Fk_#Lk4Hn5,*4n[2+n,SR
S7SSm6A52>R=RksF0k_L#54nHn,4*6[+2
,RSSSS75mAc=2R>FRskL0_kn#454H,n+*[cR2,
SSSSA7m5Rd2=s>RF_k0L4k#n,5H4[n*+,d2RS
SSmS7A25.RR=>s0Fk_#Lk4Hn5,*4n[2+.,SR
S7SSm4A52>R=RksF0k_L#54nHn,4*4[+2
,RSSSS75mAj=2R>FRskL0_kn#454H,n2*[,RR
RRRRRRRRRRRRRRRRRRRRRRRRR7RRQRuq=H>RMC_soU54*4[+(FR8IFM0R*4U[n+427,RQRuA=">Rj,j"
RRRRRRRRRRRRRRRRRRRRRRRRRRRRu7mq254RR=>IsbNH_0$L4k#n,5H.+*[4R2,7qmu5Rj2=I>RbHNs0L$_kn#45.H,*,[2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRu7mA254RR=>ssbNH_0$L4k#n,5H.+*[4R2,7Amu5Rj2=s>RbHNs0L$_kn#45.H,*2[2;R
RRRRRRRRRRRRRRFRsks0_C4o5U2*[RR<=s0Fk_#Lk4Hn5,*4n[I2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRksF0C_soU54*4[+2=R<RksF0k_L#54nHn,4*4[+2ERIC5MRs0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRs0Fk_osC5*4U[2+.RR<=s0Fk_#Lk4Hn5,*4n[2+.RCIEMsR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRsRRF_k0s5Co4[U*+Rd2<s=RF_k0L4k#n,5H4[n*+Rd2IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRFRsks0_C4o5U+*[c<2R=FRskL0_kn#454H,n+*[cI2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRksF0C_soU54*6[+2=R<RksF0k_L#54nHn,4*6[+2ERIC5MRs0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRs0Fk_osC5*4U[2+nRR<=s0Fk_#Lk4Hn5,*4n[2+nRCIEMsR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRsRRF_k0s5Co4[U*+R(2<s=RF_k0L4k#n,5H4[n*+R(2IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRFRsks0_C4o5U+*[U<2R=FRskL0_kn#454H,n+*[UI2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRksF0C_soU54*g[+2=R<RksF0k_L#54nHn,4*g[+2ERIC5MRs0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRs0Fk_osC5*4U[j+42=R<RksF0k_L#54nHn,4*4[+jI2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRksF0C_soU54*4[+4<2R=FRskL0_kn#454H,n+*[4R42IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRFRsks0_C4o5U+*[4R.2<s=RF_k0L4k#n,5H4[n*+24.RCIEMsR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRsRRF_k0s5Co4[U*+24dRR<=s0Fk_#Lk4Hn5,*4n[d+42ERIC5MRs0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRs0Fk_osC5*4U[c+42=R<RksF0k_L#54nHn,4*4[+cI2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRksF0C_soU54*4[+6<2R=FRskL0_kn#454H,n+*[4R62IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRFRsks0_C4o5U+*[4Rn2<s=RbHNs0L$_kn#45.H,*R[2IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRFRsks0_C4o5U+*[4R(2<s=RbHNs0L$_kn#45.H,*4[+2ERIC5MRs0Fk_5CMH=2RR''42DRC#'CRZ
';
RRRRRRRRRRRRRRRRkIF0C_soU54*R[2<I=RF_k0L4k#n,5H4[n*2ERIC5MRI0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRI0Fk_osC5*4U[2+4RR<=I0Fk_#Lk4Hn5,*4n[2+4RCIEMIR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRIRRF_k0s5Co4[U*+R.2<I=RF_k0L4k#n,5H4[n*+R.2IMECRF5IkC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRFRIks0_C4o5U+*[d<2R=FRIkL0_kn#454H,n+*[dI2RERCM5kIF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRkIF0C_soU54*c[+2=R<RkIF0k_L#54nHn,4*c[+2ERIC5MRI0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRI0Fk_osC5*4U[2+6RR<=I0Fk_#Lk4Hn5,*4n[2+6RCIEMIR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRIRRF_k0s5Co4[U*+Rn2<I=RF_k0L4k#n,5H4[n*+Rn2IMECRF5IkC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRFRIks0_C4o5U+*[(<2R=FRIkL0_kn#454H,n+*[(I2RERCM5kIF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRkIF0C_soU54*U[+2=R<RkIF0k_L#54nHn,4*U[+2ERIC5MRI0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRI0Fk_osC5*4U[2+gRR<=I0Fk_#Lk4Hn5,*4n[2+gRCIEMIR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRIRRF_k0s5Co4[U*+24jRR<=I0Fk_#Lk4Hn5,*4n[j+42ERIC5MRI0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRI0Fk_osC5*4U[4+42=R<RkIF0k_L#54nHn,4*4[+4I2RERCM5kIF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRkIF0C_soU54*4[+.<2R=FRIkL0_kn#454H,n+*[4R.2IMECRF5IkC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRFRIks0_C4o5U+*[4Rd2<I=RF_k0L4k#n,5H4[n*+24dRCIEMIR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRIRRF_k0s5Co4[U*+24cRR<=I0Fk_#Lk4Hn5,*4n[c+42ERIC5MRI0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRI0Fk_osC5*4U[6+42=R<RkIF0k_L#54nHn,4*4[+6I2RERCM5kIF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRkIF0C_soU54*4[+n<2R=bRIN0sH$k_L#54nH*,.[I2RERCM5kIF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRkIF0C_soU54*4[+(<2R=bRIN0sH$k_L#54nH*,.[2+4RCIEMIR5F_k0CHM52RR='24'R#CDCZR''
;
RRRRRRRRS8CMRMoCC0sNCcRz.R;
RRRRS8CMRMoCC0sNCdRzgR;
RCRRMo8RCsMCNR0Cz;dU
R
SR-RR-CRtMNCs00CRE)CRqOvRC#DDR8NMRD#CCRO0DHFoOFRVsqR)vnA4_n1d_n1d
dSzU:NRRRHV5FOEH_OCI0H8ERR=dRn2oCCMsCN0
OSzE:	RRRHV58N8s8IH0>ERRRg2oCCMsCN0
RSRRORkD:	RRFbsO#C#5iBp2S
SRoLCHSM
SHRRVBR5pCi'P0CMR8NMRiBpR'=R4R'20MEC
RSSRsRR_8N8sC_so85N8HsI8-0E4FR8IFM0RRg2<)=Rq)7758N8s8IH04E-RI8FMR0Fg
2;SRSRCRM8H
V;SMSC8sRbF#OC#ORkD
	;SRRRCRM8oCCMsCN0REzO	S;
RRRRzNdgRV:RFHsRRRHM5b8C0ME_kOl_C#DDR4-R2FR8IFM0RojRCsMCN
0CSR--Q5VRNs88I0H8ERR>gM2RCRC80OFRs0CNCsRIHR0CCLMNDNCRMF8Rkk0b0MRCNCLDRD#CCRO0DHFoOS
SSjzcNRR:H5VRNs88I0H8ERR>go2RCsMCN
0CSR--VRHGVRFsODNDRU4dUR(,#CCDOF0RVsR0HN#00MCRFL0RCoHMRosCHC#0s
C8SSSSs0Fk_5CMH<2R=4R''ERIC5MRs8_N8ss_CNo58I8sHE80-84RF0IMF2RgRH=R2DRC#'CRj
';SSSSI0Fk_5CMH<2R=4R''ERIC5MRI_N8s5CoNs88I0H8ER-48MFI0gFR2RR=HRR2CCD#R''j;S
SSsSI0M_C5RH2<W=R ERIC5MRI_N8s5CoNs88I0H8ER-48MFI0gFR2RR=HC2RDR#C';j'
SSSCRM8oCCMsCN0RjzcNS;
-Q-RVNR58I8sHE80RR<=gM2RFsRIHR0CCLMNDFCRskRF00bkRNCMLRDC#CCDOD0RFOoHRCMC8
C8SzSScR4N:VRHR85N8HsI8R0E<g=R2CRoMNCs0SC
SsSSF_k0CHM52=R<R''4;S
SSFSIkC0_M25HRR<=';4'
SSSS0Is_5CMH<2R= RW;S
SS8CMRMoCC0sNCcRz4
N;SR--tCCMsCN0RC0ERv)qRDOCDN#RM08Rs#H-0CN0#S
SS.zcNRR:VRFs[MRHRH5I8_0EM_klODCD#RR-482RF0IMFRRjoCCMsCN0
RRRRRRRRRRRRRRRR0N0skHL0\CR3lsN_VFV#\C0RRFVAv)q_.64X7d.RD:RNDLCRRH#";W"
RRRRRRRRRRRRRRRRoLCHSM
SASS)_qv6X4.dR.7:qR)vnA4_n1d_n1d
RRRRRRRRRRRRRRRRRRRRsbF0NRlb7R5Q=qR>MRH_osC5*dn[4+dRI8FMR0Fd[n*2q,R7q7)RR=>D_FII8N8sR5U8MFI0jFR27,RQ=AR>jR"jjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj,7Rq7R)A=D>RFsI_Ns8858URF0IMF2Rj,S
SShS q>R=R''4,1R1)=qR>jR''W,R =qR>sRI0M_C5,H2RiBpq>R=RiBp,hR A>R=R''4,1R1)=AR>jR''W,R =AR>jR''B,RpRiA=B>Rp
i,SSSS75mqdR42=I>RF_k0Ldk#.,5Hd[.*+2d4,SR
S7SSmdq5j=2R>FRIkL0_k.#d5dH,.+*[d,j2
SSSSq7m52.gRR=>I0Fk_#LkdH.5,*d.[g+.2
,RSSSS75mq.RU2=I>RF_k0Ldk#.,5Hd[.*+2.U,SR
S7SSm.q5(=2R>FRIkL0_k.#d5dH,.+*[.,(2
SSSSq7m52.nRR=>I0Fk_#LkdH.5,*d.[n+.2
,RSSSS75mq.R62=I>RF_k0Ldk#.,5Hd[.*+2.6,SR
S7SSm.q5c=2R>FRIkL0_k.#d5dH,.+*[.,c2
SSSSq7m52.dRR=>I0Fk_#LkdH.5,*d.[d+.2
,RSSSS75mq.R.2=I>RF_k0Ldk#.,5Hd[.*+2..,SR
S7SSm.q54=2R>FRIkL0_k.#d5dH,.+*[.,42
SSSSq7m52.jRR=>I0Fk_#LkdH.5,*d.[j+.2
,RSSSS75mq4Rg2=I>RF_k0Ldk#.,5Hd[.*+24g,SR
S7SSm4q5U=2R>FRIkL0_k.#d5dH,.+*[4,U2
SSSSq7m524(RR=>I0Fk_#LkdH.5,*d.[(+42
,RSSSS75mq4Rn2=I>RF_k0Ldk#.,5Hd[.*+24n,SR
S7SSm4q56=2R>FRIkL0_k.#d5dH,.+*[4,62
SSSSq7m524cRR=>I0Fk_#LkdH.5,*d.[c+42
,RSSSS75mq4Rd2=I>RF_k0Ldk#.,5Hd[.*+24d,SR
S7SSm4q5.=2R>FRIkL0_k.#d5dH,.+*[4,.2
SSSSq7m5244RR=>I0Fk_#LkdH.5,*d.[4+42
,RSSSS75mq4Rj2=I>RF_k0Ldk#.,5Hd[.*+24j,SR
S7SSmgq52>R=RkIF0k_L#5d.H.,d*g[+2S,
S7SSmUq52>R=RkIF0k_L#5d.H.,d*U[+2
,RSSSS75mq(=2R>FRIkL0_k.#d5dH,.+*[(R2,
SSSSq7m5Rn2=I>RF_k0Ldk#.,5Hd[.*+,n2
SSSSq7m5R62=I>RF_k0Ldk#.,5Hd[.*+,62RS
SSmS7q25cRR=>I0Fk_#LkdH.5,*d.[2+c,SR
S7SSmdq52>R=RkIF0k_L#5d.H.,d*d[+2S,
S7SSm.q52>R=RkIF0k_L#5d.H.,d*.[+2
,RSSSS75mq4=2R>FRIkL0_k.#d5dH,.+*[4R2,
SSSSq7m5Rj2=I>RF_k0Ldk#.,5Hd[.*2S,
S7SSmdA54=2R>FRskL0_k.#d5dH,.+*[d,42RS
SSmS7Aj5d2>R=RksF0k_L#5d.H.,d*d[+j
2,SSSS75mA.Rg2=s>RF_k0Ldk#.,5Hd[.*+2.g,SR
S7SSm.A5U=2R>FRskL0_k.#d5dH,.+*[.,U2RS
SSmS7A(5.2>R=RksF0k_L#5d.H.,d*.[+(
2,SSSS75mA.Rn2=s>RF_k0Ldk#.,5Hd[.*+2.n,SR
S7SSm.A56=2R>FRskL0_k.#d5dH,.+*[.,62RS
SSmS7Ac5.2>R=RksF0k_L#5d.H.,d*.[+c
2,SSSS75mA.Rd2=s>RF_k0Ldk#.,5Hd[.*+2.d,SR
S7SSm.A5.=2R>FRskL0_k.#d5dH,.+*[.,.2RS
SSmS7A45.2>R=RksF0k_L#5d.H.,d*.[+4
2,SSSS75mA.Rj2=s>RF_k0Ldk#.,5Hd[.*+2.j,SR
S7SSm4A5g=2R>FRskL0_k.#d5dH,.+*[4,g2RS
SSmS7AU542>R=RksF0k_L#5d.H.,d*4[+U
2,SSSS75mA4R(2=s>RF_k0Ldk#.,5Hd[.*+24(,SR
S7SSm4A5n=2R>FRskL0_k.#d5dH,.+*[4,n2RS
SSmS7A6542>R=RksF0k_L#5d.H.,d*4[+6
2,SSSS75mA4Rc2=s>RF_k0Ldk#.,5Hd[.*+24c,SR
S7SSm4A5d=2R>FRskL0_k.#d5dH,.+*[4,d2RS
SSmS7A.542>R=RksF0k_L#5d.H.,d*4[+.
2,SSSS75mA4R42=s>RF_k0Ldk#.,5Hd[.*+244,SR
S7SSm4A5j=2R>FRskL0_k.#d5dH,.+*[4,j2RS
SSmS7A25gRR=>s0Fk_#LkdH.5,*d.[2+g,S
SSmS7A25URR=>s0Fk_#LkdH.5,*d.[2+U,SR
S7SSm(A52>R=RksF0k_L#5d.H.,d*([+2
,RSSSS75mAn=2R>FRskL0_k.#d5dH,.+*[n
2,SSSS75mA6=2R>FRskL0_k.#d5dH,.+*[6R2,
SSSSA7m5Rc2=s>RF_k0Ldk#.,5Hd[.*+,c2RS
SSmS7A25dRR=>s0Fk_#LkdH.5,*d.[2+d,S
SSmS7A25.RR=>s0Fk_#LkdH.5,*d.[2+.,SR
S7SSm4A52>R=RksF0k_L#5d.H.,d*4[+2
,RSSSS75mAj=2R>FRskL0_k.#d5dH,.2*[,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRR7qQuRR=>HsM_Cdo5n+*[d86RF0IMFnRd*d[+.R2,7AQuRR=>"jjjj
",RRRRRRRRRRRRRRRRRRRRRRRRRRRRRmR7udq52>R=RNIbs$H0_#LkdH.5,[c*+,d2Ru7mq25.RR=>IsbNH_0$Ldk#.,5Hc+*[.
2,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRmR7u4q52>R=RNIbs$H0_#LkdH.5,[c*+,42Ru7mq25jRR=>IsbNH_0$Ldk#.,5Hc2*[,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRR7Amu5Rd2=s>RbHNs0L$_k.#d5cH,*d[+27,Rm5uA.=2R>bRsN0sH$k_L#5d.H*,c[2+.,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRR7Amu5R42=s>RbHNs0L$_k.#d5cH,*4[+27,Rm5uAj=2R>bRsN0sH$k_L#5d.H*,c[;22
RRRRRRRRRRRRRRRRsRRF_k0s5Cod[n*2=R<RksF0k_L#5d.H.,d*R[2IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRs0Fk_osC5*dn[2+4RR<=s0Fk_#LkdH.5,*d.[2+4RCIEMsR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRksF0C_son5d*.[+2=R<RksF0k_L#5d.H.,d*.[+2ERIC5MRs0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRFRsks0_Cdo5n+*[d<2R=FRskL0_k.#d5dH,.+*[dI2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRsRRF_k0s5Cod[n*+Rc2<s=RF_k0Ldk#.,5Hd[.*+Rc2IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRs0Fk_osC5*dn[2+6RR<=s0Fk_#LkdH.5,*d.[2+6RCIEMsR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRksF0C_son5d*n[+2=R<RksF0k_L#5d.H.,d*n[+2ERIC5MRs0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRFRsks0_Cdo5n+*[(<2R=FRskL0_k.#d5dH,.+*[(I2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRsRRF_k0s5Cod[n*+RU2<s=RF_k0Ldk#.,5Hd[.*+RU2IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRs0Fk_osC5*dn[2+gRR<=s0Fk_#LkdH.5,*d.[2+gRCIEMsR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRksF0C_son5d*4[+j<2R=FRskL0_k.#d5dH,.+*[4Rj2IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRs0Fk_osC5*dn[4+42=R<RksF0k_L#5d.H.,d*4[+4I2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRsRRF_k0s5Cod[n*+24.RR<=s0Fk_#LkdH.5,*d.[.+42ERIC5MRs0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRFRsks0_Cdo5n+*[4Rd2<s=RF_k0Ldk#.,5Hd[.*+24dRCIEMsR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRksF0C_son5d*4[+c<2R=FRskL0_k.#d5dH,.+*[4Rc2IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRs0Fk_osC5*dn[6+42=R<RksF0k_L#5d.H.,d*4[+6I2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRsRRF_k0s5Cod[n*+24nRR<=s0Fk_#LkdH.5,*d.[n+42ERIC5MRs0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRFRsks0_Cdo5n+*[4R(2<s=RF_k0Ldk#.,5Hd[.*+24(RCIEMsR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRksF0C_son5d*4[+U<2R=FRskL0_k.#d5dH,.+*[4RU2IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRs0Fk_osC5*dn[g+42=R<RksF0k_L#5d.H.,d*4[+gI2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRsRRF_k0s5Cod[n*+2.jRR<=s0Fk_#LkdH.5,*d.[j+.2ERIC5MRs0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRFRsks0_Cdo5n+*[.R42<s=RF_k0Ldk#.,5Hd[.*+2.4RCIEMsR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRksF0C_son5d*.[+.<2R=FRskL0_k.#d5dH,.+*[.R.2IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRs0Fk_osC5*dn[d+.2=R<RksF0k_L#5d.H.,d*.[+dI2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRsRRF_k0s5Cod[n*+2.cRR<=s0Fk_#LkdH.5,*d.[c+.2ERIC5MRs0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRFRsks0_Cdo5n+*[.R62<s=RF_k0Ldk#.,5Hd[.*+2.6RCIEMsR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRksF0C_son5d*.[+n<2R=FRskL0_k.#d5dH,.+*[.Rn2IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRs0Fk_osC5*dn[(+.2=R<RksF0k_L#5d.H.,d*.[+(I2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRsRRF_k0s5Cod[n*+2.URR<=s0Fk_#LkdH.5,*d.[U+.2ERIC5MRs0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRFRsks0_Cdo5n+*[.Rg2<s=RF_k0Ldk#.,5Hd[.*+2.gRCIEMsR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRksF0C_son5d*d[+j<2R=FRskL0_k.#d5dH,.+*[dRj2IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRs0Fk_osC5*dn[4+d2=R<RksF0k_L#5d.H.,d*d[+4I2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRsRRF_k0s5Cod[n*+2d.RR<=ssbNH_0$Ldk#.,5Hc2*[RCIEMsR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRksF0C_son5d*d[+d<2R=bRsN0sH$k_L#5d.H*,c[2+4RCIEMsR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRksF0C_son5d*d[+c<2R=bRsN0sH$k_L#5d.H*,c[2+.RCIEMsR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRksF0C_son5d*d[+6<2R=bRsN0sH$k_L#5d.H*,c[2+dRCIEMsR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRR
RRRRRRRRRRRRRRRRRI0Fk_osC5*dn[<2R=FRIkL0_k.#d5dH,.2*[RCIEMIR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRkIF0C_son5d*4[+2=R<RkIF0k_L#5d.H.,d*4[+2ERIC5MRI0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRFRIks0_Cdo5n+*[.<2R=FRIkL0_k.#d5dH,.+*[.I2RERCM5kIF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRIRRF_k0s5Cod[n*+Rd2<I=RF_k0Ldk#.,5Hd[.*+Rd2IMECRF5IkC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRI0Fk_osC5*dn[2+cRR<=I0Fk_#LkdH.5,*d.[2+cRCIEMIR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRkIF0C_son5d*6[+2=R<RkIF0k_L#5d.H.,d*6[+2ERIC5MRI0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRFRIks0_Cdo5n+*[n<2R=FRIkL0_k.#d5dH,.+*[nI2RERCM5kIF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRIRRF_k0s5Cod[n*+R(2<I=RF_k0Ldk#.,5Hd[.*+R(2IMECRF5IkC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRI0Fk_osC5*dn[2+URR<=I0Fk_#LkdH.5,*d.[2+URCIEMIR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRkIF0C_son5d*g[+2=R<RkIF0k_L#5d.H.,d*g[+2ERIC5MRI0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRFRIks0_Cdo5n+*[4Rj2<I=RF_k0Ldk#.,5Hd[.*+24jRCIEMIR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRkIF0C_son5d*4[+4<2R=FRIkL0_k.#d5dH,.+*[4R42IMECRF5IkC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRI0Fk_osC5*dn[.+42=R<RkIF0k_L#5d.H.,d*4[+.I2RERCM5kIF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRIRRF_k0s5Cod[n*+24dRR<=I0Fk_#LkdH.5,*d.[d+42ERIC5MRI0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRFRIks0_Cdo5n+*[4Rc2<I=RF_k0Ldk#.,5Hd[.*+24cRCIEMIR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRkIF0C_son5d*4[+6<2R=FRIkL0_k.#d5dH,.+*[4R62IMECRF5IkC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRI0Fk_osC5*dn[n+42=R<RkIF0k_L#5d.H.,d*4[+nI2RERCM5kIF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRIRRF_k0s5Cod[n*+24(RR<=I0Fk_#LkdH.5,*d.[(+42ERIC5MRI0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRFRIks0_Cdo5n+*[4RU2<I=RF_k0Ldk#.,5Hd[.*+24URCIEMIR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRkIF0C_son5d*4[+g<2R=FRIkL0_k.#d5dH,.+*[4Rg2IMECRF5IkC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRI0Fk_osC5*dn[j+.2=R<RkIF0k_L#5d.H.,d*.[+jI2RERCM5kIF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRIRRF_k0s5Cod[n*+2.4RR<=I0Fk_#LkdH.5,*d.[4+.2ERIC5MRI0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRFRIks0_Cdo5n+*[.R.2<I=RF_k0Ldk#.,5Hd[.*+2..RCIEMIR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRkIF0C_son5d*.[+d<2R=FRIkL0_k.#d5dH,.+*[.Rd2IMECRF5IkC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRI0Fk_osC5*dn[c+.2=R<RkIF0k_L#5d.H.,d*.[+cI2RERCM5kIF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRIRRF_k0s5Cod[n*+2.6RR<=I0Fk_#LkdH.5,*d.[6+.2ERIC5MRI0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRFRIks0_Cdo5n+*[.Rn2<I=RF_k0Ldk#.,5Hd[.*+2.nRCIEMIR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRkIF0C_son5d*.[+(<2R=FRIkL0_k.#d5dH,.+*[.R(2IMECRF5IkC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRI0Fk_osC5*dn[U+.2=R<RkIF0k_L#5d.H.,d*.[+UI2RERCM5kIF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRIRRF_k0s5Cod[n*+2.gRR<=I0Fk_#LkdH.5,*d.[g+.2ERIC5MRI0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRFRIks0_Cdo5n+*[dRj2<I=RF_k0Ldk#.,5Hd[.*+2djRCIEMIR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRkIF0C_son5d*d[+4<2R=FRIkL0_k.#d5dH,.+*[dR42IMECRF5IkC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRI0Fk_osC5*dn[.+d2=R<RNIbs$H0_#LkdH.5,[c*2ERIC5MRI0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRFRIks0_Cdo5n+*[dRd2<I=RbHNs0L$_k.#d5cH,*4[+2ERIC5MRI0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRFRIks0_Cdo5n+*[dRc2<I=RbHNs0L$_k.#d5cH,*.[+2ERIC5MRI0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRFRIks0_Cdo5n+*[dR62<I=RbHNs0L$_k.#d5cH,*d[+2ERIC5MRI0Fk_5CMH=2RR''42DRC#'CRZ
';
SSSCRM8oCCMsCN0R.zcNS;
S8CMRMoCC0sNCdRzg
N;S8CMRMoCC0sNCdRzU
N;RMRC8CRoMNCs0zCRc
d;
zRRc:cRRRHV50MFR8sN8ss_CRo2oCCMsCN0RR--oCCMsCN0RD#CCRO0s
NlRRRR-Q-RV8RN8HsI8R0E<RR6NH##o'MRj0'RFMRkk8#CR0LH#R
RRjRzRRR:H5VRNs88I0H8ERR=4o2RCsMCN
0CRRRRRRRRD_FIs8N8sR_#<"=Rjjjjj&"RR8sN_osC_j#52R;
RRRRRDRRFII_Ns88_<#R=jR"jjjj"RR&I_N8s_Co#25j;R
RRMRC8CRoMNCs0zCRjR;
RzRR4:RRRRHV58N8s8IH0=ERRR.2oCCMsCN0
RRRRRRRRIDF_8sN8#s_RR<="jjjj&"RR8sN_osC_4#5RI8FMR0Fj
2;RRRRRRRRD_FII8N8sR_#<"=Rjjjj"RR&I_N8s_Co#R548MFI0jFR2R;
RCRRMo8RCsMCNR0Cz
4;RRRRzR.R:VRHR85N8HsI8R0E=2RdRMoCC0sNCR
RRRRRRFRDIN_s8_8s#=R<Rj"jj&"RR8sN_osC_.#5RI8FMR0Fj
2;RRRRRRRRD_FII8N8sR_#<"=Rj"jjRI&RNs8_C#o_58.RF0IMF2Rj;R
RRMRC8CRoMNCs0zCR.R;
RzRRd:RRRRHV58N8s8IH0=ERRRc2oCCMsCN0
RRRRRRRRIDF_8sN8#s_RR<=""jjRs&RNs8_C#o_58dRF0IMF2Rj;R
RRRRRRFRDIN_I8_8s#=R<Rj"j"RR&I_N8s_Co#R5d8MFI0jFR2R;
RCRRMo8RCsMCNR0Cz
d;SSzc:VRHR85N8HsI8R0E=2R6RMoCC0sNCS
SD_FIs8N8sR_#<'=Rj&'RR8sN_osC_c#5RI8FMR0Fj
2;SFSDIN_I8_8s#=R<R''jRI&RNs8_C#o_58cRF0IMF2Rj;C
SMo8RCsMCNR0Cz
c;RRRRzR6R:VRHR85N8HsI8R0E>2R6RMoCC0sNCR
RRRRRRFRDIN_s8_8s#=R<R8sN_osC_6#5RI8FMR0Fj
2;RRRRRRRRD_FII8N8sR_#<I=RNs8_C#o_586RF0IMF2Rj;R
RRMRC8CRoMNCs0zCR6
;
RRRR-Q-RV8R5HsM_CRo2sHCo#s0CRh7QRHk#MBoRpRi
RzRRn:RRRRHV5M8H_osC2CRoMNCs0RC
RRRRRbRRsCFO#5#RB,piRh7Q2CRLo
HMRRRRRRRRRRRRH5VRBRpi=4R''MRN8pRBiP'CC2M0RC0EMR
RRRRRRRRRRRRRRMRH_osC_<#R=QR7hR;
RRRRRRRRRCRRMH8RVR;
RRRRRCRRMb8RsCFO#
#;RRRRCRM8oCCMsCN0R;zn
RRRRRz(RH:RVMR5F80RHsM_CRo2oCCMsCN0
RRRRRRRRRRRR_HMs_Co#=R<Rh7Q;R
RRMRC8CRoMNCs0zCR(
;
RRRR-Q-RVsR580Fk_osC2CRso0H#C7sRmRzakM#HoBRmpRi
RzRRURsR:VRHR85sF_k0s2CoRMoCC0sNCR
RRRRRRsRbF#OC#)R5_pmBis,RF_k0s_Co#L2RCMoH
RRRRRRRRRRRRRHV5m)_BRpi=4R''MRN8_R)miBp'CCPMR020MEC
RRRRRRRRRRRRRRRR7)_mRza<s=RF_k0s_Co#R;
RRRRRRRRRCRRMH8RVR;
RRRRRCRRMb8RsCFO#
#;RRRRCRM8oCCMsCN0RszU;R
RRgRzs:RRRRHV50MFRFs8ks0_CRo2oCCMsCN0
RRRRRRRRRRRR7)_mRza<s=RF_k0s_Co#R;
RCRRMo8RCsMCNR0Cz;gs
z
SURIR:VRHR85IF_k0s2CoRMoCC0sNCR
RRRRRRsRbF#OC#WR5_pmBiI,RF_k0s_Co#L2RCMoH
RRRRRRRRRRRRRHV5mW_BRpi=4R''MRN8_RWmiBp'CCPMR020MEC
RRRRRRRRRRRRRRRR7W_mRza<I=RF_k0s_Co#R;
RRRRRRRRRCRRMH8RVR;
RRRRRCRRMb8RsCFO#
#;RRRRCRM8oCCMsCN0RIzU;R
RRgRzI:RRRRHV50MFRFI8ks0_CRo2oCCMsCN0
RRRRRRRRRRRR7W_mRza<I=RF_k0s_Co#R;
RCRRMo8RCsMCNR0Cz;gI
R
RR-R-RRQV58sN8ss_CRo2sHCo#s0CR7q7)#RkHRMoB
piRRRRzR4jRH:RVsR5Ns88_osC2CRoMNCs0RC
RRRRRbRRsCFO#5#R)B_mpRi,)7q7)L2RCMoH
RRRRRRRRRRRRRHV5m)_BRpi=4R''MRN8_R)miBp'CCPMR020MEC
RRRRRRRRRRRRRRRR8sN_osC_<#R=qR)757)Ns88I0H8ER-48MFI0jFR2R;
RRRRRRRRRCRRMH8RVR;
RRRRRCRRMb8RsCFO#
#;RRRRCRM8oCCMsCN0Rjz4;R
RR4Rz4RR:H5VRMRF0s8N8sC_soo2RCsMCN
0CRRRRRRRRRRRRs_N8s_Co#=R<R7)q7
);RRRRCRM8oCCMsCN0R4z4;R

R-RR-VRQRN5I8_8ss2CoRosCHC#0s7Rq7k)R#oHMRiBp
RRRR.z4RRR:H5VRI8N8sC_soo2RCsMCN
0CRRRRRRRRbOsFCR##5iBp,qRW727)RoLCHRM
RRRRRRRRRHRRVBR5p=iRR''4R8NMRiBp'CCPMR020MEC
RRRRRRRRRRRRRRRR8IN_osC_<#R=qRW757)Ns88I0H8ER-48MFI0jFR2R;
RRRRRRRRRCRRMH8RVR;
RRRRRCRRMb8RsCFO#
#;RRRRCRM8oCCMsCN0R.z4;R
RR4RzdRR:H5VRMRF0I8N8sC_soo2RCsMCN
0CRRRRRRRRRRRRI_N8s_Co#=R<R7Wq7
);RRRRCRM8oCCMsCN0Rdz4;R
RRRRRRRR
R-RR-CRtMNCs00CRE)CRqOvRC#DDR8NMRD#CCRO0DHFoOR
RR4RzcRR:VRFsHMRHRk5MlC_ODnD_cRR-482RF0IMFRRjoCCMsCN0
RRRRR--Q5VRNs88I0H8ERR>6M2RCRC80OFRs0CNCsRIHR0CCLMNDNCRMF8Rkk0b0MRCNCLDRD#CCRO0DHFoOR
RRRRRR4Rz6RR:H5VRNs88I0H8ERR>no2RCsMCN
0CRRRRRRRRRRRRRRRRs0Fk__CM#25HRR<='R4'IMECRN5s8C_so5_#Ns88I0H8ER-48MFI0nFR2RR=HC2RDR#C';j'
SSSSkIF0M_C_H#52=R<R''4RCIEMIR5Ns8_C#o_58N8s8IH04E-RI8FMR0Fn=2RRRH2CCD#R''j;R
RRRRRRRRRRRRRRsRI0M_C_H#52=R<RRW IMECRN5I8C_so5_#Ns88I0H8ER-48MFI0nFR2RR=HC2RDR#C';j'
RRRRRRRR8CMRMoCC0sNC4Rz6R;
R-RR-VRQR85N8HsI8R0E<6=R2FRMRHIs0CCRMDNLCsRFR0FkbRk0CLMND#CRCODC0FRDoRHOM8CCCR8
RRRRRzRR4:nRRRHV58N8s8IH0<ER=2RnRMoCC0sNCR
RRRRRRRRRRRRRRFRskC0_M5_#H<2R=4R''S;
SISSF_k0C#M_5RH2<'=R4
';RRRRRRRRRRRRRRRRI_s0C#M_5RH2<W=R R;
RRRRRCRRMo8RCsMCNR0Cz;4n
RRRRR--tCCMsCN0RC0ERv)qRDOCDN#RM08Rs#H-0CN0#R
RRRRRR4Rz(RR:VRFs[MRHRH5I8R0E-2R4RI8FMR0FjCRoMNCs0RC
RRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)RzqcvnRD:RNDLCRRH#"a17"RR&HCM0o'CsHolNCH5I820ER"&R7&"RR0HMCsoC'NHloHC5*2ncR"&RW&"RR0HMCsoC'NHlo[C52RR&"R "&MRH0CCosl'HN5oCo_C0C_M880CbEH55+*42nRc,80CbER22&XR""RR&HCM0o'CsHolNC+5[4
2;RRRRRRRRRRRRLHCoMR
RRRRRRRRRR)RzqcvnRX:R)nqvc7X4RR
RRRRRRRRRRRRRRFRbsl0RN5bR7>R=R_HMs_Co#25[,jRqRR=>D_FII8N8s5_#jR2,q=4R>FRDIN_I8_8s#254,.RqRR=>D_FII8N8s5_#.
2,RRRRRRRRRRRRRRRRRRRRRRRRRdRqRR=>D_FII8N8s5_#dR2,q=cR>FRDIN_I8_8s#25c,6RqRR=>D_FII8N8s5_#6R2,
SSSSRSSR)7uq=jR>FRDIN_s8_8s#25j,uR7)Rq4=D>RFsI_Ns88_4#527,Ru.)qRR=>D_FIs8N8s5_#.
2,SSSSSRSR7qu)d>R=RIDF_8sN8#s_5,d2R)7uq=cR>FRDIN_s8_8s#25c,uR7)Rq6=D>RFsI_Ns88_6#52
,RSSSSSRSRW= R>sRI0M_C_H#52W,RBRpi=B>RpRi,7Rum=s>RF_k0L_k#n5c#H2,[,uR1m>R=RkIF0k_L#c_n#,5H[;22
RRRRRRRRRRRRRRRRksF0C_so5_#[<2R=FRskL0_kn#_cH#5,R[2IMECRF5skC0_M5_#H=2RR''42DRC#'CRZ
';SSSSI0Fk_osC_[#52=R<RkIF0k_L#c_n#,5H[I2RERCM5kIF0M_C_H#52RR='24'R#CDCZR''R;
RRRRRCRRMo8RCsMCNR0Cz;4(
RRRRMRC8CRoMNCs0zCR4Rc;RRRRRRRRR
RRRRRRRRR
R-RR-CRtMNCs0NCRRRd.I8FsRC8CbqR)vCRODHDRVbRNbbsFs0HNCRRRRRRRRRRRRRRR
RRRRUz4RH:RVMR5kOl_C_DDd=.RRR42oCCMsCN0
RRRRR--Q5VRNs88I0H8ERR>(M2RCRC80OFRs0CNCsRIHR0CCLMNDNCRMF8Rkk0b0MRCNCLDRD#CCRO0DHFoOR
RRRRRR4Rzg:NRRRHV58N8s8IH0>ERRRn2oCCMsCN0
RRRRRRRRRRRRRRRRksF0M_C_Rd.<'=R4I'RERCM5N5s8C_so5_#Ns88I0H8ER-48MFI0nFR2RR=M_klODCD_2ncR8NMRN5s8C_so5_#6=2RR''j2C2RDR#C';j'
SSSSkIF0M_C_Rd.<'=R4I'RERCM5N5I8C_so5_#Ns88I0H8ER-48MFI0nFR2RR=M_klODCD_2ncR8NMRN5I8C_so5_#6=2RR''j2C2RDR#C';j'
RRRRRRRRRRRRRRRR0Is__CMd<.R= RWRCIEM5R5I_N8s_Co#85N8HsI8-0E4FR8IFM0RRn2=kRMlC_ODnD_cN2RM58RI_N8s_Co#256R'=Rj2'2R#CDCjR''R;
RRRRRCRRMo8RCsMCNR0CzN4g;R
RRRRRR4Rzg:LRRRHV58N8s8IH0=ERRNnRMM8RkOl_C_DDn=cRRRj2oCCMsCN0
RRRRRRRRRRRRRRRRksF0M_C_Rd.<'=R4I'RERCM5N5s8C_so5_#6=2RR''j2C2RDR#C';j'
SSSSkIF0M_C_Rd.<'=R4I'RERCM5N5I8C_so5_#6=2RR''j2C2RDR#C';j'
RRRRRRRRRRRRRRRR0Is__CMd<.R= RWRCIEM5R5I_N8s_Co#256R'=Rj2'2R#CDCjR''R;
RRRRRCRRMo8RCsMCNR0CzL4g;RRRRR--Q5VRNs88I0H8E=R<RR62MIFRsCH0RNCMLRDCFFsRkk0b0MRCNCLDRD#CCRO0DHFoOCRMC88C
RRRRRRRRjz.RH:RVNR58I8sHE80RR<=6o2RCsMCN
0CRRRRRRRRRRRRRRRRs0Fk__CMd<.R=4R''S;
SISSF_k0CdM_.=R<R''4;R
RRRRRRRRRRRRRRsRI0M_C_Rd.<W=R R;
RRRRRCRRMo8RCsMCNR0Cz;.j
RRRRR--tCCMsCN0RC0ERv)qRDOCDMRN8sR0H0-#N
0CRRRRRRRRzR.4:FRVsRR[H5MRI0H8ERR-482RF0IMFRRjoCCMsCN0
RRRRRRRRRRRR0N0skHL0\CR3lsN_VFV#\C0RRFVzv)qd:.RRLDNCHDR#1R"7Ra"&MRH0CCosl'HN5oCI0H8E&2RR""7RH&RMo0CCHs'lCNo5lMk_DOCDc_n*2ncR"&RW&"RR0HMCsoC'NHlo[C52RR&"R "&MRH0CCosl'HN5oCo_C0C_M880CbEk5MlC_ODnD_cc*nRd+R.8,RCEb02&2RR""XRH&RMo0CCHs'lCNo54[+2R;
RRRRRRRRRLRRCMoH
RRRRRRRRRRRRqz)vRd.:)RXq.vdXR47
RRRRRRRRRRRRRRRRsbF0NRlb7R5RR=>HsM_C#o_5,[2RRqj=D>RFII_Ns88_j#52q,R4>R=RIDF_8IN8#s_5,42RRq.=D>RFII_Ns88_.#52R,
RRRRRRRRRRRRRRRRRRRRRRRRRRqd=D>RFII_Ns88_d#52q,Rc>R=RIDF_8IN8#s_5,c2RS
SSSSSRuR7)Rqj=D>RFsI_Ns88_j#527,Ru4)qRR=>D_FIs8N8s5_#4R2,7qu).>R=RIDF_8sN8#s_5,.2
SSSSRSSR)7uq=dR>FRDIN_s8_8s#25d,uR7)Rqc=D>RFsI_Ns88_c#52
,RSSSSSRSRW= R>sRI0M_C_,d.RpWBi>R=RiBp,uR7m>R=RksF0k_L#._d#k5MlC_ODdD_.2,[,uR1m>R=RkIF0k_L#._d#k5MlC_ODdD_.2,[2R;
RRRRRRRRRRRRRsRRF_k0s_Co#25[RR<=s0Fk_#Lk_#d.5lMk_DOCD._d,R[2IMECRF5skC0_M._dR'=R4R'2CCD#R''Z;S
SSFSIks0_C#o_5R[2<I=RF_k0L_k#d5.#M_klODCD_,d.[I2RERCM5kIF0M_C_Rd.=4R''C2RDR#C';Z'
RRRRRRRRMRC8CRoMNCs0zCR.
4;RRRRR8CMRMoCC0sNC4RzUR;RRRRRRRRR
R
RR-R-RMtCC0sNCRRN4InRFRs88bCCRv)qRDOCDVRHRbNbssFbHCN0RRRRRRRRRRRRR
RRRRRRzR..:VRHRk5MlC_OD4D_nRR=4o2RCsMCN
0CRRRR-Q-RVNR58I8sHE80R6>R2CRMC08RFsROCCN0RHIs0CCRMDNLCMRN8kRF00bkRNCMLRDC#CCDOD0RFOoH
RRRRRRRRdz.NRR:H5VRNs88I0H8ERR>nMRN8kRMlC_ODdD_.RR=4o2RCsMCN
0CRRRRRRRRRRRRRRRRs0Fk__CM4<nR=4R''ERIC5MR58sN_osC_N#58I8sHE80-84RF0IMF2RnRM=RkOl_C_DDnRc2NRM858sN_osC_6#52RR='24'R8NMRN5s8C_so5_#c=2RR''j2C2RDR#C';j'
SSSSkIF0M_C_R4n<'=R4I'RERCM5N5I8C_so5_#Ns88I0H8ER-48MFI0nFR2RR=M_klODCD_2ncR8NMRN5I8C_so5_#6=2RR''42MRN8IR5Ns8_C#o_5Rc2=jR''R22CCD#R''j;R
RRRRRRRRRRRRRRsRI0M_C_R4n<W=R ERIC5MR58IN_osC_N#58I8sHE80-84RF0IMF2RnRM=RkOl_C_DDnRc2NRM858IN_osC_6#52RR='24'R8NMRN5I8C_so5_#c=2RR''j2C2RDR#C';j'
RRRRRRRR8CMRMoCC0sNC.Rzd
N;RRRRRRRRzL.dRH:RVNR58I8sHE80Rn>RR8NMRlMk_DOCD._dRR/=4o2RCsMCN
0CRRRRRRRRRRRRRRRRs0Fk__CM4<nR=4R''ERIC5MR58sN_osC_N#58I8sHE80-84RF0IMF2RnRM=RkOl_C_DDnRc2NRM858sN_osC_6#52RR='2j'R8NMRN5s8C_so5_#c=2RR''j2C2RDR#C';j'
SSSSkIF0M_C_R4n<'=R4I'RERCM5N5I8C_so5_#Ns88I0H8ER-48MFI0nFR2RR=M_klODCD_2ncR8NMRN5I8C_so5_#6=2RR''j2MRN8IR5Ns8_C#o_5Rc2=jR''R22CCD#R''j;R
RRRRRRRRRRRRRRsRI0M_C_R4n<W=R ERIC5MR58IN_osC_N#58I8sHE80-84RF0IMF2RnRM=RkOl_C_DDnRc2NRM858IN_osC_6#52RR='2j'R8NMRN5I8C_so5_#c=2RR''j2C2RDR#C';j'
RRRRRRRR8CMRMoCC0sNC.Rzd
L;RRRRRRRRzO.dRH:RVNR58I8sHE80Rn=RR8NMRlMk_DOCD._dR4=R2CRoMNCs0RC
RRRRRRRRRRRRRsRRF_k0C4M_n=R<R''4RCIEM5R5s_N8s_Co#256R'=R4R'2NRM858sN_osC_c#52RR='2j'2DRC#'CRj
';SSSSI0Fk__CM4<nR=4R''ERIC5MR58IN_osC_6#52RR='24'R8NMRN5I8C_so5_#c=2RR''j2C2RDR#C';j'
RRRRRRRRRRRRRRRR0Is__CM4<nR= RWRCIEM5R5I_N8s_Co#256R'=R4R'2NRM858IN_osC_c#52RR='2j'2DRC#'CRj
';RRRRRRRRCRM8oCCMsCN0Rdz.OR;
RRRRRzRR.Rd8:VRHR85N8HsI8R0E=RR6NRM8M_klODCD_Rd./4=R2CRoMNCs0RC
RRRRRRRRRRRRRsRRF_k0C4M_n=R<R''4RCIEM5R5s_N8s_Co#85N8HsI8-0E4FR8IFM0RRc2=kRMlC_ODdD_.R22CCD#R''j;S
SSFSIkC0_Mn_4RR<='R4'IMECRI55Ns8_C#o_58N8s8IH04E-RI8FMR0Fc=2RRlMk_DOCD._d2C2RDR#C';j'
RRRRRRRRRRRRRRRR0Is__CM4<nR= RWRCIEM5R5I_N8s_Co#85N8HsI8-0E4FR8IFM0RRc2=kRMlC_ODdD_.R22CCD#R''j;R
RRRRRRMRC8CRoMNCs0zCR.;d8RRRR-Q-RVNR58I8sHE80RR<=6M2RFsRIHR0CCLMNDFCRskRF00bkRNCMLRDC#CCDOD0RFOoHRCMC8
C8RRRRRRRRzR.c:VRHR85N8HsI8R0E<c=R2CRoMNCs0RC
RRRRRRRRRRRRRsRRF_k0C4M_n=R<R''4;S
SSFSIkC0_Mn_4RR<=';4'
RRRRRRRRRRRRRRRR0Is__CM4<nR= RW;R
RRRRRRMRC8CRoMNCs0zCR.
c;RRRR-t-RCsMCNR0C0REC)RqvODCDR8NMRH0s-N#00RC
RRRRRzRR.:6RRsVFRH[RMIR5HE80R4-R2FR8IFM0RojRCsMCN
0CRRRRRRRRRRRRNs00H0LkC3R\s_NlF#VVCR0\FzVR)4qvnRR:DCNLD#RHR7"1a&"RR0HMCsoC'NHloIC5HE802RR&"R7"&MRH0CCosl'HN5oCM_klODCD_*ncn+cRRlMk_DOCD._d*2d.R"&RW&"RR0HMCsoC'NHlo[C52RR&"R "&MRH0CCosl'HN5oCo_C0C_M880CbEk5MlC_ODnD_cc*nRM+RkOl_C_DDdd.*.RR+4Rn,80CbER22&XR""RR&HCM0o'CsHolNC+5[4
2;RRRRRRRRRRRRLHCoMR
RRRRRRRRRR)Rzqnv4R):Rqnv4XR47
RRRRRRRRRRRRRRRRsbF0NRlb7R5RR=>HsM_C#o_5,[2RRqj=D>RFII_Ns88_j#52q,R4>R=RIDF_8IN8#s_5,42RRq.=D>RFII_Ns88_.#52R,
RRRRRRRRRRRRRRRRRRRRRRRRRRqd=D>RFII_Ns88_d#527,Ruj)qRR=>D_FIs8N8s5_#jR2,7qu)4>R=RIDF_8sN8#s_5,42R)7uq=.R>FRDIN_s8_8s#25.,S
SSSSSRuR7)Rqd=D>RFsI_Ns88_d#52W,R >R=R0Is__CM4Rn,WiBpRR=>B,piRm7uRR=>s0Fk_#Lk_#4n5lMk_DOCDn_4,,[2Rm1uRR=>I0Fk_#Lk_#4n5lMk_DOCDn_4,2[2;R
RRRRRRRRRRRRRRFRsks0_C#o_5R[2<s=RF_k0L_k#45n#M_klODCD_,4n[I2RERCM5ksF0M_C_R4n=4R''C2RDR#C';Z'
SSSSkIF0C_so5_#[<2R=FRIkL0_k4#_nM#5kOl_C_DD4[n,2ERIC5MRI0Fk__CM4=nRR''42DRC#'CRZ
';RRRRRRRRCRM8oCCMsCN0R6z.;R
RRMRC8CRoMNCs0zCR.R.;R
RRRMRC8CRoMNCs0zCRc
c;CRM8NEsOHO0C0CksR_MFsOI_E	CO;-

--
----
-R--p0N#RbHlDCClM00NHRFMH8#RCkVND-0
-R--#CCDOs0_NNl
sHOE00COkRsC#CCDOs0_NFlRVqR)vW_)uR_)HV#
k0MOHRFMo_C0C_M880CbEH5#x:CRR0HMCsoCR8;RCEb0RH:RMo0CCRs2skC0sHMRMo0CCHsR#N
PsLHNDlCRH#M_HRxC:MRH0CCos=R:R
j;LHCoMR
Rl_HM#CHxRR:=80CbER;
RRHV5x#HCRR<80CbE02RE
CMRRRRl_HM#CHxRR:=#CHx;R
RCRM8H
V;RCRs0MksRMlH_x#HCC;
Mo8RCC0_M88_CEb0;F
OMN#0MM0RkOl_C#DDRH:RMo0CC:sR=5R580CbERR-442/nR2;RRRRRRRRR-RR-RRyF)VRqnv4XR47ODCD#CRMC88C
b0$CkRF0k_L#$_0bHCR#sRNsRN$5lMk_DOCD8#RF0IMF,RjR8IH04E-RI8FMR0FjF2RV0R#8F_Do;HO
o#HMRNDs0Fk_#LkRF:RkL0_k0#_$;bCRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RR.7NNss$VRFR8s_FRk05bHMk00RFsR0H0-#N#0C2H
#oDMNRksF0M_CR#:R0D8_FOoH_OPC05FsM_klODCD#FR8IFM0R;j2RRRRR-RR-MRCNCLD#FRVssR0H0-#N#0C
o#HMRNDI0Fk_RCM:0R#8F_Do_HOP0COFMs5kOl_C#DDRI8FMR0Fj
2;#MHoNIDRF_k0LRk#:kRF0k_L#$_0bRC;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--.N7Rs$sNRRFVIF_8k50RHkMb0FR0RH0s-N#002C#
o#HMRNDI_s0C:MRR8#0_oDFHPO_CFO0sk5MlC_ODRD#8MFI0jFR2R;RRRRRR-R-RHIs0CCRMDNLCV#RFCsRNROEsRFIF)VRqOvRC#DD
o#HMRNDHsM_C:oRR8#0_oDFHPO_CFO0sH5I8-0E4FR8IFM0R;j2RRRRRRRRR-R-RCk#8FR0RosCHC#0sQR7h#R
HNoMDFRsks0_C:oRR8#0_oDFHPO_CFO0sH5I8-0E4FR8IFM0R;j2RRRRRRRR-k-R#RC80sFRC#oH0RCs)m_7z#a
HNoMDFRIks0_C:oRR8#0_oDFHPO_CFO0sH5I8-0E4FR8IFM0R;j2RRRRRRRR-k-R#RC80sFRC#oH0RCsWm_7z#a
HNoMDNRs8C_soRR:#_08DHFoOC_POs0F58N8s8IH04E-RI8FMR0FjR2;RRRR-k-R#RC80sFRC#oH0RCs)7q7)H
#oDMNR8IN_osCR#:R0D8_FOoH_OPC05FsNs88I0H8ER-48MFI0jFR2R;RR-RR-#RkC08RFCRso0H#CWsRq)77
o#HMRNDD_FIs8N8sRR:#_08DHFoOC_POs0F58dRF0IMF2Rj;RRRRRRRRRRRR-R-R8sN8LsRHR0#HkMb0FR0Rv)qRDOCD5#RcHRL0s#RCHJks2C8
o#HMRNDD_FII8N8sRR:#_08DHFoOC_POs0F58dRF0IMF2Rj;RRRRRRRRRRRR-R-R8IN8LsRHR0#HkMb0FR0Rv)qRDOCD5#RcHRL0s#RCHJks2C8
0N0skHL0\CR3lsN_VFV#\C0R#:R0MsHo
;
LHCoMR

R-RR-VRQR8N8s8IH0<ERRNcR#o#HMjR''FR0RkkM#RC8L#H0
RRRRRz4RH:RVNR58I8sHE80R4=R2CRoMNCs0RC
RRRRRDRRFsI_Ns88RR<="jjj"RR&s_N8s5Coj
2;RRRRRRRRD_FII8N8s=R<Rj"jj&"RR8IN_osC5;j2
RRRR8CMRMoCC0sNC4Rz;R
RR.RzRRR:H5VRNs88I0H8ERR=.o2RCsMCN
0CRRRRRRRRD_FIs8N8s=R<Rj"j"RR&s_N8s5Co4FR8IFM0R;j2
RRRRRRRRIDF_8IN8<sR=jR"j&"RR8IN_osC584RF0IMF2Rj;R
RRMRC8CRoMNCs0zCR.R;
RzRRd:RRRRHV58N8s8IH0=ERRRd2oCCMsCN0
RRRRRRRRIDF_8sN8<sR=jR''RR&s_N8s5Co.FR8IFM0R;j2
RRRRRRRRIDF_8IN8<sR=jR''RR&I_N8s5Co.FR8IFM0R;j2
RRRR8CMRMoCC0sNCdRz;R
RRcRzRRR:H5VRNs88I0H8ERR>do2RCsMCN
0CRRRRRRRRD_FIs8N8s=R<R8sN_osC58dRF0IMF2Rj;R
RRRRRRFRDIN_I8R8s<I=RNs8_Cdo5RI8FMR0Fj
2;RRRRCRM8oCCMsCN0R;zc
R
RR-R-RRQV5M8H_osC2CRso0H#C7sRQkhR#oHMRiBp
RRRRRz6RH:RV8R5HsM_CRo2oCCMsCN0
RRRRRRRRFbsO#C#Rp5Bi7,RQRh2LHCoMR
RRRRRRRRRRVRHRp5BiRR='R4'NRM8B'piCMPC002RE
CMRRRRRRRRRRRRRRRRHsM_C<oR=QR7hR;
RRRRRRRRRCRRMH8RVR;
RRRRRCRRMb8RsCFO#
#;RRRRCRM8oCCMsCN0R;z6
RRRRRznRH:RVMR5F80RHsM_CRo2oCCMsCN0
RRRRRRRRRRRR_HMsRCo<7=RQ
h;RRRRCRM8oCCMsCN0R;zn
R
RR-R-RRQV5ksF0C_sos2RC#oH0RCs7amzRHk#MmoRB
piRRRRzR(sRH:RVsR580Fk_osC2CRoMNCs0RC
RRRRRbRRsCFO#5#R)B_mpRi,s0Fk_osC2CRLo
HMRRRRRRRRRRRRH5VR)B_mp=iRR''4R8NMRm)_B'piCMPC002RE
CMRRRRRRRRRRRRRRRR)m_7z<aR=FRsks0_C
o;RRRRRRRRRRRRCRM8H
V;RRRRRRRRCRM8bOsFC;##
RRRR8CMRMoCC0sNC(RzsR;
RzRRURsR:VRHRF5M08RsF_k0s2CoRMoCC0sNCR
RRRRRRRRRR_R)7amzRR<=s0Fk_osC;R
RRMRC8CRoMNCs0zCRU
s;
RRRRR--Q5VRs0Fk_osC2CRso0H#C7sRmRzakM#HoBRmpRi
RzRR(RIR:VRHR85IF_k0s2CoRMoCC0sNCR
RRRRRRsRbF#OC#WR5_pmBiI,RF_k0s2CoRoLCHRM
RRRRRRRRRHRRVWR5_pmBiRR='R4'NRM8WB_mpCi'P0CM2ER0CRM
RRRRRRRRRRRRRWRR_z7ma=R<RkIF0C_soR;
RRRRRRRRRCRRMH8RVR;
RRRRRCRRMb8RsCFO#
#;RRRRCRM8oCCMsCN0RIz(;R
RRURzI:RRRRHV50MFRFI8ks0_CRo2oCCMsCN0
RRRRRRRRRRRR7W_mRza<I=RF_k0s;Co
RRRR8CMRMoCC0sNCURzI
;
RRRR-Q-RVsR5Ns88_osC2CRso0H#C)sRq)77RHk#MmoRB
piRRRRzRgR:VRHRN5s8_8ss2CoRMoCC0sNCR
RRRRRRsRbF#OC#)R5_pmBi),Rq)772CRLo
HMRRRRRRRRRRRRH5VR)B_mp=iRR''4R8NMRm)_B'piCMPC002RE
CMRRRRRRRRRRRRRRRRs_N8sRCo<)=Rq)7758N8s8IH04E-RI8FMR0Fj
2;RRRRRRRRRRRRCRM8H
V;RRRRRRRRCRM8bOsFC;##
RRRR8CMRMoCC0sNCgRz;R
RR4RzjRR:H5VRMRF0s8N8sC_soo2RCsMCN
0CRRRRRRRRRRRRs_N8sRCo<)=Rq)77;R
RRMRC8CRoMNCs0zCR4
j;RRRRRRRR
RRRRR--Q5VRI8N8sC_sos2RC#oH0RCsW7q7)#RkHRMoB
piRRRRzR46RH:RVIR5Ns88_osC2CRoMNCs0RC
RRRRRbRRsCFO#5#RB,piR7Wq7R)2LHCoMR
RRRRRRRRRRVRHRp5BiRR='R4'NRM8B'piCMPC002RE
CMRRRRRRRRRRRRRRRRI_N8sRCo<W=Rq)7758N8s8IH04E-RI8FMR0Fj
2;RRRRRRRRRRRRCRM8H
V;RRRRRRRRCRM8bOsFC;##
RRRR8CMRMoCC0sNC4Rz6R;
RzRR4:nRRRHV50MFR8IN8ss_CRo2oCCMsCN0
RRRRRRRRRRRR8IN_osCRR<=W7q7)R;
RCRRMo8RCsMCNR0Cz;4n
R
RR-R-RMtCC0sNCER0CqR)vCRODRD#NRM8#CCDOD0RFOoH
RRRR4z4RV:RFHsRRRHMM_klODCD#FR8IFM0RojRCsMCN
0CRRRRRRRR-Q-RVNR58I8sHE80Rc>R2CRMC08RFsROCCN0RHIs0CCRMDNLCMRN8kRF00bkRNCMLRDC#CCDOD0RFOoH
RRRRRRRR.z4RH:RVNR58I8sHE80Rc>R2CRoMNCs0RC
RRRRRRRRRRRRRsRRF_k0CHM52=R<R''4RCIEMsR5Ns8_CNo58I8sHE80-84RF0IMF2RcRH=R2DRC#'CRj
';RRRRRRRRRRRRRRRRI0Fk_5CMH<2R=4R''ERIC5MRI_N8s5CoNs88I0H8ER-48MFI0cFR2RR=HC2RDR#C';j'
RRRRRRRRRRRRRRRR0Is_5CMH<2R= RWRCIEMIR5Ns8_CNo58I8sHE80-84RF0IMF2RcRH=R2DRC#'CRj
';RRRRRRRRCRM8oCCMsCN0R.z4;R
RRRRRR-R-RRQV58N8s8IH0<ER=2RcRRMFI0sHCMRCNCLDRRFsFbk0kC0RMDNLCCR#D0CORoDFHMORCCC88R
RRRRRR4RzdRR:H5VRNs88I0H8E=R<RRc2oCCMsCN0
RRRRRRRRRRRRRRRRksF0M_C5RH2<'=R4
';RRRRRRRRRRRRRRRRI0Fk_5CMH<2R=4R''R;
RRRRRRRRRRRRRIRRsC0_M25HRR<=W
 ;RRRRRRRRRRRRCRM8oCCMsCN0Rdz4;R
RR-R-RCtMsCN0RC0ERv)qRDOCDN#RM08Rs#H-0CN0#R
RRRRRR4RzcRR:VRFs[MRHRH5I8R0E-2R4RI8FMR0FjCRoMNCs0RC
RRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)Rzq:vRRLDNCHDR#1R"7Ra"&MRH0CCosl'HN5oCI0H8E&2RR""7RH&RMo0CCHs'lCNo54H*n&2RR""WRH&RMo0CCHs'lCNo5R[2& R""RR&HCM0o'CsHolNCC5o0M_C8C_8b50E54H+2n*4,CR8b20E2RR&"RX"&MRH0CCosl'HN5oC[2+4;R
RRRRRRRRRRCRLo
HMRRRRRRRRRRRRzv)q:qR)vX4n4
7RRRRRRRRRRRRRRRRRb0FsRblNRR57=H>RMC_so25[,jRqRR=>D_FII8N8s25j,4RqRR=>D_FII8N8s254,.RqRR=>D_FII8N8s25.,R
RRRRRRRRRRRRRRRRRRRRRRRRRq=dR>FRDIN_I858sdR2,7qu)j>R=RIDF_8sN8js527,Ru4)qRR=>D_FIs8N8s254,RR
RRRRRRRRRRRRRRRRRRRRRRRRR)7uq=.R>FRDIN_s858s.R2,7qu)d>R=RIDF_8sN8ds52W,R >R=R0Is_5CMHR2,
RRRRRRRRRRRRRRRRRRRRRRRRWRRBRpi=B>RpRi,7Rum=s>RF_k0L5k#H2,[,uR1m>R=RkIF0k_L#,5H[;22
RRRRRRRRRRRRksF0C_so25[RR<=s0Fk_#Lk5[H,2ERIC5MRs0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRI0Fk_osC5R[2<I=RF_k0L5k#H2,[RCIEMIR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRCRRMo8RCsMCNR0Cz;4c
RRRRRRRR8CMRMoCC0sNC4Rz4R;
RRRRRRRRRRRRRRRRRRRRRRRRRRRR
8CMRONsECH0Os0kCCR#D0CO_lsN;



