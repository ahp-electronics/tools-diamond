library verilog;
use verilog.vl_types.all;
entity cfg_register is
    port(
        fsd_persistn_progn: out    vl_logic;
        fsd_persist_initn: out    vl_logic;
        fsd_persist_done: out    vl_logic;
        fsd_persistn_jtag: out    vl_logic;
        fsd_persistn_sspi: out    vl_logic;
        fsd_persistn_i2c: out    vl_logic;
        fsd_persist_mspi: out    vl_logic;
        fsd_boot_sel    : out    vl_logic_vector(2 downto 0);
        sd_i2c_addr     : out    vl_logic_vector(7 downto 0);
        sd_i2c_deg      : out    vl_logic;
        sd_i2c_deg_sel  : out    vl_logic;
        sd_dec_only     : out    vl_logic;
        sd_pwd_ufm      : out    vl_logic;
        sd_pwd_en       : out    vl_logic;
        sd_pwd_all      : out    vl_logic;
        sd_cid_en       : out    vl_logic;
        sd_vrbp_en      : out    vl_logic;
        sd_pwd_mismatch : out    vl_logic;
        sd_trim0        : out    vl_logic_vector(127 downto 0);
        sd_trim1        : out    vl_logic_vector(127 downto 0);
        ctrl0           : out    vl_logic_vector(31 downto 0);
        ctrl1           : out    vl_logic_vector(31 downto 0);
        dryrun_spi_flash_addr: out    vl_logic_vector(23 downto 0);
        cidcode         : out    vl_logic_vector(31 downto 0);
        uidcode         : out    vl_logic_vector(63 downto 0);
        ctrl_m_addr2    : out    vl_logic_vector(23 downto 0);
        comp_dic        : out    vl_logic_vector(127 downto 0);
        key_byte        : out    vl_logic_vector(7 downto 0);
        sd_aes_key      : out    vl_logic_vector(255 downto 0);
        sd_auth_en      : out    vl_logic_vector(1 downto 0);
        sd_rand_noise   : out    vl_logic;
        sd_rand_aes     : out    vl_logic;
        sd_secplus_cfg0 : out    vl_logic;
        sd_done_cfg0    : out    vl_logic;
        sd_authdone_cfg0: out    vl_logic;
        sd_ues_cfg0     : out    vl_logic_vector(31 downto 0);
        sd_secplus_cfg1 : out    vl_logic;
        sd_done_cfg1    : out    vl_logic;
        sd_authdone_cfg1: out    vl_logic;
        sd_ues_cfg1     : out    vl_logic_vector(31 downto 0);
        sd_sec_read_sram: out    vl_logic;
        sd_sec_erase_sram: out    vl_logic;
        sd_sec_read_cfg0: out    vl_logic;
        sd_sec_prog_cfg0: out    vl_logic;
        sd_sec_erase_cfg0: out    vl_logic;
        sd_sec_read_cfg1: out    vl_logic;
        sd_sec_prog_cfg1: out    vl_logic;
        sd_sec_erase_cfg1: out    vl_logic;
        sd_sec_read_fea : out    vl_logic;
        sd_sec_prog_fea : out    vl_logic;
        sd_sec_erase_fea: out    vl_logic;
        sd_sec_read_trim: out    vl_logic;
        sd_sec_prog_trim: out    vl_logic;
        sd_sec_erase_trim: out    vl_logic;
        sd_sec_read_pubkey: out    vl_logic;
        sd_sec_prog_pubkey: out    vl_logic;
        sd_sec_erase_pubkey: out    vl_logic;
        sd_sec_read_aeskey: out    vl_logic;
        sd_sec_prog_aeskey: out    vl_logic;
        sd_sec_erase_aeskey: out    vl_logic;
        sd_sec_read_csec: out    vl_logic;
        sd_sec_prog_csec: out    vl_logic;
        sd_sec_erase_csec: out    vl_logic;
        sd_sec_read_usec: out    vl_logic;
        sd_sec_prog_usec: out    vl_logic;
        sd_sec_erase_usec: out    vl_logic;
        sd_sec_read_ufm0: out    vl_logic;
        sd_sec_prog_ufm0: out    vl_logic;
        sd_sec_erase_ufm0: out    vl_logic;
        sd_sec_read_ufm1: out    vl_logic;
        sd_sec_prog_ufm1: out    vl_logic;
        sd_sec_erase_ufm1: out    vl_logic;
        sd_sec_read_ufm2: out    vl_logic;
        sd_sec_prog_ufm2: out    vl_logic;
        sd_sec_erase_ufm2: out    vl_logic;
        sd_sec_read_ufm3: out    vl_logic;
        sd_sec_prog_ufm3: out    vl_logic;
        sd_sec_erase_ufm3: out    vl_logic;
        sd_sec_hlock_cfg0: out    vl_logic;
        sd_sec_hlock_cfg1: out    vl_logic;
        sd_sec_hlock_trim: out    vl_logic;
        sd_sec_hlock_fea: out    vl_logic;
        sd_sec_hlock_pubkey: out    vl_logic;
        sd_sec_hlock_aeskey: out    vl_logic;
        sd_sec_hlock_csec: out    vl_logic;
        sd_sec_hlock_ufm0: out    vl_logic;
        sd_sec_hlock_ufm1: out    vl_logic;
        sd_sec_hlock_ufm2: out    vl_logic;
        sd_sec_hlock_ufm3: out    vl_logic;
        sd_sec_hlock_usec: out    vl_logic;
        sd_sec_hlock_sram: out    vl_logic;
        sd_sec_hlock_jtag: out    vl_logic;
        sd_sec_jtag     : out    vl_logic_vector(1 downto 0);
        sd_sec_hlock_sspi: out    vl_logic;
        sd_sec_sspi     : out    vl_logic_vector(1 downto 0);
        sd_sec_hlock_si2c: out    vl_logic;
        sd_sec_si2c     : out    vl_logic_vector(1 downto 0);
        sd_sec_hlock_bspi: out    vl_logic;
        sd_sec_bspi     : out    vl_logic;
        sd_sec_hlock_bi2c: out    vl_logic;
        sd_sec_bi2c     : out    vl_logic;
        mt_freq_cnt     : out    vl_logic_vector(15 downto 0);
        cfg_reg_dat     : out    vl_logic_vector(127 downto 0);
        id_err          : out    vl_logic;
        njs_invalid_err : out    vl_logic;
        buf128_dat      : out    vl_logic_vector(127 downto 0);
        cfg_i2c_dat     : out    vl_logic_vector(15 downto 0);
        cfg_ctrl0_upd   : out    vl_logic;
        cfg0_latter     : out    vl_logic;
        dryrun_ues      : out    vl_logic_vector(31 downto 0);
        sd_ues          : out    vl_logic_vector(31 downto 0);
        sd_done         : out    vl_logic;
        sec_read_alt_sram: out    vl_logic;
        sec_prog_alt_sram: out    vl_logic;
        sd_uds_trn      : out    vl_logic_vector(127 downto 0);
        uds_trn_blank   : out    vl_logic;
        hse_trn_valid   : out    vl_logic;
        sec_ucode_set   : out    vl_logic_vector(31 downto 0);
        pwdMismatchAtCheck: out    vl_logic;
        por             : in     vl_logic;
        por_sec         : in     vl_logic;
        por_trim        : in     vl_logic;
        smclk           : in     vl_logic;
        smclk_scan_off  : in     vl_logic;
        nj_rst_flag     : in     vl_logic;
        scanen          : in     vl_logic;
        CTRL0_DEFAULT   : in     vl_logic_vector(31 downto 0);
        CTRL1_DEFAULT   : in     vl_logic_vector(31 downto 0);
        finish_cdm      : in     vl_logic;
        fl_start_cdm    : in     vl_logic;
        ASSP_EN         : in     vl_logic;
        ENC_ONLY_EN     : in     vl_logic;
        p_slave         : in     vl_logic;
        bg_cmp_out      : in     vl_logic;
        proc_ring_osc   : in     vl_logic;
        mfg_freq_sel    : in     vl_logic;
        mfg_bkgrndft_en : in     vl_logic;
        buf128_int      : in     vl_logic_vector(127 downto 0);
        contxt_dat      : in     vl_logic_vector(7 downto 0);
        nj_exec_b       : in     vl_logic;
        isc_exec_e      : in     vl_logic;
        idcode_err      : in     vl_logic;
        bse_active      : in     vl_logic;
        mfg_en          : in     vl_logic;
        access_sudo     : in     vl_logic;
        access_safe     : in     vl_logic;
        rti_r           : in     vl_logic;
        upir_ss_r       : in     vl_logic;
        exit1dr_ss_r    : in     vl_logic;
        ref_start       : in     vl_logic;
        nj_rst_ctrl01   : in     vl_logic;
        rst_ctrl01_onfail: in     vl_logic;
        bse_err_rst     : in     vl_logic;
        fl_udss0_authdone_qual: in     vl_logic;
        fl_udss1_authdone_qual: in     vl_logic;
        lsc_prog_uds_qual: in     vl_logic;
        dryrun_prog_ucode_qual: in     vl_logic;
        dryrun_check_exec: in     vl_logic;
        access_flash_manu: in     vl_logic;
        current_sector  : in     vl_logic_vector(11 downto 0);
        fl_load_trim0   : in     vl_logic;
        fl_load_trim1   : in     vl_logic;
        fl_load_pes     : in     vl_logic;
        fl_load_mes     : in     vl_logic;
        fl_load_pwd     : in     vl_logic;
        fl_load_fea     : in     vl_logic;
        fl_load_feabits : in     vl_logic;
        fl_load_udss0   : in     vl_logic;
        fl_load_ufs0    : in     vl_logic;
        fl_load_tss     : in     vl_logic;
        fl_load_fss     : in     vl_logic;
        fl_load_uds_trn : in     vl_logic;
        fl_erase_cfg0   : in     vl_logic;
        fl_erase_ufm0   : in     vl_logic;
        fl_erase_trim   : in     vl_logic;
        fl_erase_fea    : in     vl_logic;
        fl_load_pkey0   : in     vl_logic;
        fl_load_pkey1   : in     vl_logic;
        fl_load_pkey2   : in     vl_logic;
        fl_load_pkey3   : in     vl_logic;
        fl_load_udss1   : in     vl_logic;
        fl_load_ufs1    : in     vl_logic;
        fl_load_pks     : in     vl_logic;
        fl_load_css     : in     vl_logic;
        fl_load_csec    : in     vl_logic;
        fl_erase_cfg1   : in     vl_logic;
        fl_erase_ufm1   : in     vl_logic;
        fl_erase_pubkey : in     vl_logic;
        fl_erase_csec   : in     vl_logic;
        fl_load_akey0   : in     vl_logic;
        fl_load_akey1   : in     vl_logic;
        fl_load_ufs2    : in     vl_logic;
        fl_load_ufs3    : in     vl_logic;
        fl_load_aks     : in     vl_logic;
        fl_load_uss     : in     vl_logic;
        fl_load_usec    : in     vl_logic;
        fl_erase_ufm2   : in     vl_logic;
        fl_erase_ufm3   : in     vl_logic;
        fl_erase_aeskey : in     vl_logic;
        fl_erase_usec   : in     vl_logic;
        verify_id_qual  : in     vl_logic;
        lsc_prog_ctrl0_qual: in     vl_logic;
        lsc_prog_ctrl1_qual: in     vl_logic;
        prog_dryrun_addr_qual: in     vl_logic;
        lsc_write_comp_dic_qual: in     vl_logic;
        lsc_shift_password_qual: in     vl_logic;
        isc_prog_done_qual: in     vl_logic;
        isc_prog_sec_qual: in     vl_logic;
        isc_prog_secplus_qual: in     vl_logic;
        isc_prog_ucode_qual: in     vl_logic;
        lsc_prog_authmode_qual: in     vl_logic;
        lsc_prog_aesfea_qual: in     vl_logic;
        lsc_prog_password_qual: in     vl_logic;
        lsc_prog_cipher_key0_qual: in     vl_logic;
        lsc_prog_cipher_key1_qual: in     vl_logic;
        lsc_prog_pubkey0_qual: in     vl_logic;
        lsc_prog_pubkey1_qual: in     vl_logic;
        lsc_prog_pubkey2_qual: in     vl_logic;
        lsc_prog_pubkey3_qual: in     vl_logic;
        lsc_prog_feature_qual: in     vl_logic;
        lsc_prog_feabits_qual: in     vl_logic;
        lsc_prog_trim0_qual: in     vl_logic;
        lsc_prog_trim1_qual: in     vl_logic;
        lsc_prog_pes_qual: in     vl_logic;
        lsc_prog_mes_qual: in     vl_logic;
        lsc_prog_csec_qual: in     vl_logic;
        lsc_prog_usec_qual: in     vl_logic;
        lsc_read_authmode_qual: in     vl_logic;
        lsc_read_aesfea_qual: in     vl_logic;
        lsc_read_password_qual: in     vl_logic;
        lsc_read_cipher_key0_qual: in     vl_logic;
        lsc_read_cipher_key1_qual: in     vl_logic;
        lsc_read_pubkey0_qual: in     vl_logic;
        lsc_read_pubkey1_qual: in     vl_logic;
        lsc_read_pubkey2_qual: in     vl_logic;
        lsc_read_pubkey3_qual: in     vl_logic;
        lsc_read_feature_qual: in     vl_logic;
        lsc_read_feabits_qual: in     vl_logic;
        lsc_read_trim0_qual: in     vl_logic;
        lsc_read_trim1_qual: in     vl_logic;
        lsc_read_pes_qual: in     vl_logic;
        lsc_read_mes_qual: in     vl_logic;
        lsc_read_usec_qual: in     vl_logic;
        lsc_read_csec_qual: in     vl_logic;
        fl_write_addr_qual: in     vl_logic;
        fl_disable_done0_qual: in     vl_logic;
        fl_disable_done1_qual: in     vl_logic;
        mfg_mdata_qual  : in     vl_logic;
        mfg_mtrim_qual  : in     vl_logic;
        cmd_altsec_ufm3 : in     vl_logic;
        cmd_altsec_ufm2 : in     vl_logic;
        cmd_altsec_ufm1 : in     vl_logic;
        cmd_altsec_ufm0 : in     vl_logic;
        cmd_altsec_jtag : in     vl_logic;
        cmd_altsec_sspi : in     vl_logic;
        cmd_altsec_si2c : in     vl_logic;
        cmd_altsec_bspi : in     vl_logic;
        cmd_altsec_bi2c : in     vl_logic;
        cmd_altsec_sram : in     vl_logic;
        cmd_altsec_cfg0 : in     vl_logic;
        cmd_altsec_cfg1 : in     vl_logic;
        cmd_altsec_pubkey: in     vl_logic;
        cmd_altsec_aeskey: in     vl_logic;
        cmd_altsec_trim : in     vl_logic;
        cmd_altsec_fea  : in     vl_logic;
        cmd_altsec_usec : in     vl_logic;
        cmd_altsec_csec : in     vl_logic;
        sed_prog_ctrl0_qual: in     vl_logic;
        sed_prog_ctrl1_qual: in     vl_logic;
        sed_write_comp_dic_qual: in     vl_logic;
        njbse_rst_flag  : in     vl_logic;
        isc_disable_exec: in     vl_logic;
        exec_buf        : in     vl_logic_vector(127 downto 0);
        key_rst_sync    : in     vl_logic;
        key_shift_en    : in     vl_logic;
        njs_invalid_c   : in     vl_logic;
        hse_trn_dat     : in     vl_logic_vector(127 downto 0)
    );
end cfg_register;
