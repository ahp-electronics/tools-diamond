-- Remove REN for MS;
-- Added arc for AS_LSB;
-- Modified the array element to pass MTI;
-- REV 1.1;
LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.VITAL_timing.all;
USE IEEE.VITAL_primitives.all;
 
 
package VLOGTOVITAL_TABLES is
 
---------------------------------------------------------------------------------
-- Local type declaration
---------------------------------------------------------------------------------

    TYPE edge_table IS ARRAY (std_ulogic, std_ulogic) OF boolean ;

---------------------------------------------------------------------------------
-- Contants Specifications
-- posedge, negedge
---------------------------------------------------------------------------------
    CONSTANT POSEDGE : edge_table := (
    --      ---------------------------------------------------------
    --      |  U      X      0      1      Z      W      L      H      - |   |
    --      ---------------------------------------------------------
            ( FALSE, FALSE, FALSE, TRUE, FALSE, FALSE, FALSE, FALSE, FALSE ), -- | U |
            ( FALSE, FALSE, FALSE, TRUE, FALSE, FALSE, FALSE, FALSE, FALSE ), -- | X |
            ( FALSE, TRUE,  FALSE, TRUE, FALSE, FALSE, FALSE, FALSE, FALSE ), -- | 0 |
            ( FALSE, FALSE, FALSE, FALSE,FALSE, FALSE, FALSE, FALSE, FALSE ), -- | 1 |
            ( FALSE, FALSE, FALSE, TRUE, FALSE, FALSE, FALSE, FALSE, FALSE ), -- | Z |
            ( FALSE, FALSE, FALSE, TRUE, FALSE, FALSE, FALSE, FALSE, FALSE ), -- | W |
            ( FALSE, TRUE,  FALSE, TRUE, FALSE, FALSE, FALSE, FALSE, FALSE ), -- | L |
            ( FALSE, FALSE, FALSE, FALSE,FALSE, FALSE, FALSE, FALSE, FALSE ), -- | H |
            ( FALSE, FALSE, FALSE, FALSE,FALSE, FALSE, FALSE, FALSE, FALSE )  -- | - |
        );

    CONSTANT NEGEDGE : edge_table := (
    --      ---------------------------------------------------- -----
    --      |  U    X    0    1    Z    W    L    H    - |   |
    --      ---------------------------------------------------- -----
            ( FALSE, FALSE, TRUE, FALSE, FALSE, FALSE, FALSE, FALSE, FALSE ), -- | U |
            ( FALSE, FALSE, TRUE, FALSE, FALSE, FALSE, FALSE, FALSE, FALSE ), -- | X |
            ( FALSE, FALSE, FALSE,FALSE, FALSE, FALSE, FALSE, FALSE, FALSE ), -- | 0 |
            ( FALSE, TRUE,  TRUE, FALSE, FALSE, FALSE, FALSE, FALSE, FALSE ), -- | 1 |
            ( FALSE, FALSE, TRUE, FALSE, FALSE, FALSE, FALSE, FALSE, FALSE ), -- | Z |
            ( FALSE, FALSE, TRUE, FALSE, FALSE, FALSE, FALSE, FALSE, FALSE ), -- | W |
            ( FALSE, FALSE, FALSE,FALSE, FALSE, FALSE, FALSE, FALSE, FALSE ), -- | L |
            ( FALSE, TRUE,  TRUE, FALSE, FALSE, FALSE, FALSE, FALSE, FALSE ), -- | H |
            ( FALSE, FALSE, FALSE,FALSE, FALSE, FALSE, FALSE, FALSE, FALSE )  -- | - |
        );

        -------------------------------------------------------------------------------
        --State Table Declaration
        -------------------------------------------------------------------------------

	CONSTANT dfftab : VitalStateTableType := (
	-- D CLK R S lstSt Q
	( '-', '-', '0', '1', '-', '0' ),
	( '-', '-', '1', '0', '-', '1' ),
	( '1', '/', '1', '-', '-', '1' ),
	( '0', '/', '-', '1', '-', '0' ),
	( '1', '-', '1', '*', '1', '1' ),
	( '-', '0', '1', '*', '1', '1' ),
	( '-', '1', '1', '*', '1', '1' ),
	( '1', '-', '0', '\', '0', 'X' ),---
	( '-', '0', '0', '\', '0', 'X' ),---
	( '-', '1', '0', '\', '0', 'X' ),---
	( '0', '-', '*', '1', '0', '0' ),
	( '-', '0', '*', '1', '0', '0' ),
	( '-', '1', '*', '1', '0', '0' ),
	( '0', '-', '\', '0', '1', 'X' ),--
	( '-', '0', '\', '0', '1', 'X' ),--
	( '-', '1', '\', '0', '1', 'X' ),--
	( '1', 'R', '1', '1', '1', '1' ),
	( '0', 'R', '1', '1', '0', '0' ),
	( '-', '\', '-', '-', '-', 'S' ),
	( '-', 'v', '-', '-', '-', 'S' ),
	( '0', 'r', '-', '-', '0', 'S' ),
	( '0', 'f', '-', '-', '0', 'S' ),
	( '1', 'r', '-', '-', '1', 'S' ),
	( '1', 'f', '-', '-', '1', 'S' ),
	( '*', '1', '-', '-', '-', 'S' ),
	( '*', '0', '-', '-', '-', 'S' ),
	( 'S', 'S', 'S', 'S', '-', 'S' ),
	( 'r', 'S', 'S', 'S', '-', 'X' ),
	( 'f', 'S', 'S', 'S', '-', 'X' ),
	( 'X', 'S', 'S', 'S', '-', 'S' ),
	( 'S', 'r', 'S', 'S', '-', 'X' ),
	( 'S', 'f', 'S', 'S', '-', 'X' ),
	( 'S', 'X', 'S', 'S', '-', 'S' ),
	( 'r', 'X', 'S', 'S', '-', 'X' ),
	( 'f', 'X', 'S', 'S', '-', 'X' ),
	( 'X', 'r', 'S', 'S', '-', 'X' ),
	( 'X', 'f', 'S', 'S', '-', 'X' ),
	( 'X', 'X', 'S', 'S', '-', 'S' ),
	( 'S', 'S', 'r', 'S', '-', 'X' ),
	( 'S', 'S', 'f', 'S', '-', 'X' ),
	( 'S', 'S', 'X', 'S', '-', 'S' ),
	( 'r', 'S', 'X', 'S', '-', 'X' ),
	( 'f', 'S', 'X', 'S', '-', 'X' ),
	( 'X', 'S', 'r', 'S', '-', 'X' ),
	( 'X', 'S', 'f', 'S', '-', 'X' ),
	( 'X', 'S', 'X', 'S', '-', 'S' ),
	( 'S', 'r', 'X', 'S', '-', 'X' ),
	( 'S', 'f', 'X', 'S', '-', 'X' ),
	( 'S', 'X', 'r', 'S', '-', 'X' ),
	( 'S', 'X', 'f', 'S', '-', 'X' ),
	( 'S', 'X', 'X', 'S', '-', 'S' ),
	( 'r', 'X', 'X', 'S', '-', 'X' ),
	( 'f', 'X', 'X', 'S', '-', 'X' ),
	( 'X', 'r', 'X', 'S', '-', 'X' ),
	( 'X', 'f', 'X', 'S', '-', 'X' ),
	( 'X', 'X', 'r', 'S', '-', 'X' ),
	( 'X', 'X', 'f', 'S', '-', 'X' ),
	( 'X', 'X', 'X', 'S', '-', 'S' ),
	( 'S', 'S', 'S', 'r', '-', 'X' ),
	( 'S', 'S', 'S', 'f', '-', 'X' ),
	( 'S', 'S', 'S', 'X', '-', 'S' ),
	( 'r', 'S', 'S', 'X', '-', 'X' ),
	( 'f', 'S', 'S', 'X', '-', 'X' ),
	( 'X', 'S', 'S', 'r', '-', 'X' ),
	( 'X', 'S', 'S', 'f', '-', 'X' ),
	( 'X', 'S', 'S', 'X', '-', 'S' ),
	( 'S', 'r', 'S', 'X', '-', 'X' ),
	( 'S', 'f', 'S', 'X', '-', 'X' ),
	( 'S', 'X', 'S', 'r', '-', 'X' ),
	( 'S', 'X', 'S', 'f', '-', 'X' ),
	( 'S', 'X', 'S', 'X', '-', 'S' ),
	( 'r', 'X', 'S', 'X', '-', 'X' ),
	( 'f', 'X', 'S', 'X', '-', 'X' ),
	( 'X', 'r', 'S', 'X', '-', 'X' ),
	( 'X', 'f', 'S', 'X', '-', 'X' ),
	( 'X', 'X', 'S', 'r', '-', 'X' ),
	( 'X', 'X', 'S', 'f', '-', 'X' ),
	( 'X', 'X', 'S', 'X', '-', 'S' ),
	( 'S', 'S', 'r', 'X', '-', 'X' ),
	( 'S', 'S', 'f', 'X', '-', 'X' ),
	( 'S', 'S', 'X', 'r', '-', 'X' ),
	( 'S', 'S', 'X', 'f', '-', 'X' ),
	( 'S', 'S', 'X', 'X', '-', 'S' ),
	( 'r', 'S', 'X', 'X', '-', 'X' ),
	( 'f', 'S', 'X', 'X', '-', 'X' ),
	( 'X', 'S', 'r', 'X', '-', 'X' ),
	( 'X', 'S', 'f', 'X', '-', 'X' ),
	( 'X', 'S', 'X', 'r', '-', 'X' ),
	( 'X', 'S', 'X', 'f', '-', 'X' ),
	( 'X', 'S', 'X', 'X', '-', 'S' ),
	( 'S', 'r', 'X', 'X', '-', 'X' ),
	( 'S', 'f', 'X', 'X', '-', 'X' ),
	( 'S', 'X', 'r', 'X', '-', 'X' ),
	( 'S', 'X', 'f', 'X', '-', 'X' ),
	( 'S', 'X', 'X', 'r', '-', 'X' ),
	( 'S', 'X', 'X', 'f', '-', 'X' ),
	( 'S', 'X', 'X', 'X', '-', 'S' ),
	( 'r', 'X', 'X', 'X', '-', 'X' ),
	( 'f', 'X', 'X', 'X', '-', 'X' ),
	( 'X', 'r', 'X', 'X', '-', 'X' ),
	( 'X', 'f', 'X', 'X', '-', 'X' ),
	( 'X', 'X', 'r', 'X', '-', 'X' ),
	( 'X', 'X', 'f', 'X', '-', 'X' ),
	( 'X', 'X', 'X', 'r', '-', 'X' ),
	( 'X', 'X', 'X', 'f', '-', 'X' ),
	( 'X', 'X', 'X', 'X', '-', 'S' ) );


	-------------------------------------------------------------------------------
	--State Table Declaration
	-------------------------------------------------------------------------------
	CONSTANT latchtab : VitalStateTableType := (
	-- D LAT R S lstSt Q
	( '-', '-', '0', '1', '-', '0' ),
	( '-', '-', '1', '0', '-', '1' ),
	( '*', '0', '1', '1', '-', 'S' ),
	( '-', '\', '1', '1', '-', 'S' ),
	( '-', 'v', '1', '1', '-', 'S' ),
	( '-', 'f', '1', '1', '-', 'S' ),
	( '0', '^', '-', '1', '-', '0' ),
	( '1', '^', '1', '-', '-', '1' ),
	( '0', 'r', '1', '1', '0', '0' ),
	( '1', 'r', '1', '1', '1', '1' ),
	( '\', '1', '-', '1', '-', '0' ),
	( 'v', '1', '-', '1', '-', '0' ),
	( '/', '1', '1', '-', '-', '1' ),
	( '^', '1', '1', '-', '-', '1' ),
	( '0', '/', '-', '1', '-', '0' ),
	( '1', '/', '1', '-', '-', '1' ),
	( '-', '0', '1', '/', '-', 'S' ),
	( '-', '0', '1', '^', '-', 'S' ),
	( '-', '0', '/', '1', '-', 'S' ),
	( '-', '0', '^', '1', '-', 'S' ),
	( '0', '1', '-', '/', '-', '0' ),
	( '0', '1', '-', '^', '-', '0' ),
	( '1', '1', '/', '-', '-', '1' ),
	( '1', '1', '^', '-', '-', '1' ),
	( '1', '1', '1', '/', '-', '1' ),
	( '1', '1', '1', '^', '-', '1' ),
	( '0', '1', '/', '1', '-', '0' ),
	( '0', '1', '^', '1', '-', '0' ),
	( '/', 'X', '1', '-', '1', '1' ),
	( '^', 'X', '1', '-', '1', '1' ),
	( '\', 'X', '-', '1', '0', '0' ),
	( 'v', 'X', '-', '1', '0', '0' ),
	( 'S', 'S', 'S', 'S', '-', 'S' ),
	( 'r', 'S', 'S', 'S', '-', 'X' ),
	( 'f', 'S', 'S', 'S', '-', 'X' ),
	( 'X', 'S', 'S', 'S', '-', 'S' ),
	( 'S', 'r', 'S', 'S', '-', 'X' ),
	( 'S', 'f', 'S', 'S', '-', 'X' ),
	( 'S', 'X', 'S', 'S', '-', 'S' ),
	( 'r', 'X', 'S', 'S', '-', 'X' ),
	( 'f', 'X', 'S', 'S', '-', 'X' ),
	( 'X', 'r', 'S', 'S', '-', 'X' ),
	( 'X', 'f', 'S', 'S', '-', 'X' ),
	( 'X', 'X', 'S', 'S', '-', 'S' ),
	( 'S', 'S', 'r', 'S', '-', 'X' ),
	( 'S', 'S', 'f', 'S', '-', 'X' ),
	( 'S', 'S', 'X', 'S', '-', 'S' ),
	( 'r', 'S', 'X', 'S', '-', 'X' ),
	( 'f', 'S', 'X', 'S', '-', 'X' ),
	( 'X', 'S', 'r', 'S', '-', 'X' ),
	( 'X', 'S', 'f', 'S', '-', 'X' ),
	( 'X', 'S', 'X', 'S', '-', 'S' ),
	( 'S', 'r', 'X', 'S', '-', 'X' ),
	( 'S', 'f', 'X', 'S', '-', 'X' ),
	( 'S', 'X', 'r', 'S', '-', 'X' ),
	( 'S', 'X', 'f', 'S', '-', 'X' ),
	( 'S', 'X', 'X', 'S', '-', 'S' ),
	( 'r', 'X', 'X', 'S', '-', 'X' ),
	( 'f', 'X', 'X', 'S', '-', 'X' ),
	( 'X', 'r', 'X', 'S', '-', 'X' ),
	( 'X', 'f', 'X', 'S', '-', 'X' ),
	( 'X', 'X', 'r', 'S', '-', 'X' ),
	( 'X', 'X', 'f', 'S', '-', 'X' ),
	( 'X', 'X', 'X', 'S', '-', 'S' ),
	( 'S', 'S', 'S', 'r', '-', 'X' ),
	( 'S', 'S', 'S', 'f', '-', 'X' ),
	( 'S', 'S', 'S', 'X', '-', 'S' ),
	( 'r', 'S', 'S', 'X', '-', 'X' ),
	( 'f', 'S', 'S', 'X', '-', 'X' ),
	( 'X', 'S', 'S', 'r', '-', 'X' ),
	( 'X', 'S', 'S', 'f', '-', 'X' ),
	( 'X', 'S', 'S', 'X', '-', 'S' ),
	( 'S', 'r', 'S', 'X', '-', 'X' ),
	( 'S', 'f', 'S', 'X', '-', 'X' ),
	( 'S', 'X', 'S', 'r', '-', 'X' ),
	( 'S', 'X', 'S', 'f', '-', 'X' ),
	( 'S', 'X', 'S', 'X', '-', 'S' ),
	( 'r', 'X', 'S', 'X', '-', 'X' ),
	( 'f', 'X', 'S', 'X', '-', 'X' ),
	( 'X', 'r', 'S', 'X', '-', 'X' ),
	( 'X', 'f', 'S', 'X', '-', 'X' ),
	( 'X', 'X', 'S', 'r', '-', 'X' ),
	( 'X', 'X', 'S', 'f', '-', 'X' ),
	( 'X', 'X', 'S', 'X', '-', 'S' ),
	( 'S', 'S', 'r', 'X', '-', 'X' ),
	( 'S', 'S', 'f', 'X', '-', 'X' ),
	( 'S', 'S', 'X', 'r', '-', 'X' ),
	( 'S', 'S', 'X', 'f', '-', 'X' ),
	( 'S', 'S', 'X', 'X', '-', 'S' ),
	( 'r', 'S', 'X', 'X', '-', 'X' ),
	( 'f', 'S', 'X', 'X', '-', 'X' ),
	( 'X', 'S', 'r', 'X', '-', 'X' ),
	( 'X', 'S', 'f', 'X', '-', 'X' ),
	( 'X', 'S', 'X', 'r', '-', 'X' ),
	( 'X', 'S', 'X', 'f', '-', 'X' ),
	( 'X', 'S', 'X', 'X', '-', 'S' ),
	( 'S', 'r', 'X', 'X', '-', 'X' ),
	( 'S', 'f', 'X', 'X', '-', 'X' ),
	( 'S', 'X', 'r', 'X', '-', 'X' ),
	( 'S', 'X', 'f', 'X', '-', 'X' ),
	( 'S', 'X', 'X', 'r', '-', 'X' ),
	( 'S', 'X', 'X', 'f', '-', 'X' ),
	( 'S', 'X', 'X', 'X', '-', 'S' ),
	( 'r', 'X', 'X', 'X', '-', 'X' ),
	( 'f', 'X', 'X', 'X', '-', 'X' ),
	( 'X', 'r', 'X', 'X', '-', 'X' ),
	( 'X', 'f', 'X', 'X', '-', 'X' ),
	( 'X', 'X', 'r', 'X', '-', 'X' ),
	( 'X', 'X', 'f', 'X', '-', 'X' ),
	( 'X', 'X', 'X', 'r', '-', 'X' ),
	( 'X', 'X', 'X', 'f', '-', 'X' ),
	( 'X', 'X', 'X', 'X', '-', 'S' ) );


	-------------------------------------------------------------------------------
	--State Table Declaration
	-------------------------------------------------------------------------------
	CONSTANT jkfftab : VitalStateTableType := (
	-- CLK J K S R lstSt Q
	( '-', '-', '-', '0', '1', '-', '1' ),
	( '-', '-', '-', '1', '0', '-', '0' ),
	( '-', '-', '-', '*', '1', '1', '1' ),
	( '-', '-', '-', '1', '*', '0', '0' ),
	( '/', '0', '0', '1', '1', '-', 'S' ),
	( '/', '0', '1', '1', '1', '-', '0' ),
	( '/', '1', '0', '1', '1', '-', '1' ),
	( '/', '1', '1', '1', '1', '1', '0' ),
	( '/', '1', '1', '1', '1', '0', '1' ),
	( '\', '-', '-', '-', '-', '-', 'S' ),
	( 'B', '*', '-', '-', '-', '-', 'S' ),
	( 'B', '-', '*', '-', '-', '-', 'S' ),
	( 'R', '0', '0', '1', '1', '-', 'S' ),
	( 'R', '0', '-', '1', '-', '0', 'S' ),
	( 'R', '-', '0', '-', '1', '1', 'S' ),
	( 'v', '-', '-', '-', '-', '-', 'S' ),
	( 'f', '0', '0', '1', '1', '-', 'S' ),
	( 'f', '0', '-', '1', '-', '0', 'S' ),
	( 'f', '-', '0', '-', '1', '1', 'S' ),
	( 'X', '*', '0', '-', '1', '1', 'S' ),
	( 'X', '0', '*', '1', '-', '0', 'S' ),
	( 'S', 'S', 'S', 'S', 'S', '-', 'S' ),
	( 'r', 'S', 'S', 'S', 'S', '-', 'X' ),
	( 'f', 'S', 'S', 'S', 'S', '-', 'X' ),
	( 'X', 'S', 'S', 'S', 'S', '-', 'S' ),
	( 'S', 'r', 'S', 'S', 'S', '-', 'X' ),
	( 'S', 'f', 'S', 'S', 'S', '-', 'X' ),
	( 'S', 'X', 'S', 'S', 'S', '-', 'S' ),
	( 'r', 'X', 'S', 'S', 'S', '-', 'X' ),
	( 'f', 'X', 'S', 'S', 'S', '-', 'X' ),
	( 'X', 'r', 'S', 'S', 'S', '-', 'X' ),
	( 'X', 'f', 'S', 'S', 'S', '-', 'X' ),
	( 'X', 'X', 'S', 'S', 'S', '-', 'S' ),
	( 'S', 'S', 'r', 'S', 'S', '-', 'X' ),
	( 'S', 'S', 'f', 'S', 'S', '-', 'X' ),
	( 'S', 'S', 'X', 'S', 'S', '-', 'S' ),
	( 'r', 'S', 'X', 'S', 'S', '-', 'X' ),
	( 'f', 'S', 'X', 'S', 'S', '-', 'X' ),
	( 'X', 'S', 'r', 'S', 'S', '-', 'X' ),
	( 'X', 'S', 'f', 'S', 'S', '-', 'X' ),
	( 'X', 'S', 'X', 'S', 'S', '-', 'S' ),
	( 'S', 'r', 'X', 'S', 'S', '-', 'X' ),
	( 'S', 'f', 'X', 'S', 'S', '-', 'X' ),
	( 'S', 'X', 'r', 'S', 'S', '-', 'X' ),
	( 'S', 'X', 'f', 'S', 'S', '-', 'X' ),
	( 'S', 'X', 'X', 'S', 'S', '-', 'S' ),
	( 'r', 'X', 'X', 'S', 'S', '-', 'X' ),
	( 'f', 'X', 'X', 'S', 'S', '-', 'X' ),
	( 'X', 'r', 'X', 'S', 'S', '-', 'X' ),
	( 'X', 'f', 'X', 'S', 'S', '-', 'X' ),
	( 'X', 'X', 'r', 'S', 'S', '-', 'X' ),
	( 'X', 'X', 'f', 'S', 'S', '-', 'X' ),
	( 'X', 'X', 'X', 'S', 'S', '-', 'S' ),
	( 'S', 'S', 'S', 'r', 'S', '-', 'X' ),
	( 'S', 'S', 'S', 'f', 'S', '-', 'X' ),
	( 'S', 'S', 'S', 'X', 'S', '-', 'S' ),
	( 'r', 'S', 'S', 'X', 'S', '-', 'X' ),
	( 'f', 'S', 'S', 'X', 'S', '-', 'X' ),
	( 'X', 'S', 'S', 'r', 'S', '-', 'X' ),
	( 'X', 'S', 'S', 'f', 'S', '-', 'X' ),
	( 'X', 'S', 'S', 'X', 'S', '-', 'S' ),
	( 'S', 'r', 'S', 'X', 'S', '-', 'X' ),
	( 'S', 'f', 'S', 'X', 'S', '-', 'X' ),
	( 'S', 'X', 'S', 'r', 'S', '-', 'X' ),
	( 'S', 'X', 'S', 'f', 'S', '-', 'X' ),
	( 'S', 'X', 'S', 'X', 'S', '-', 'S' ),
	( 'r', 'X', 'S', 'X', 'S', '-', 'X' ),
	( 'f', 'X', 'S', 'X', 'S', '-', 'X' ),
	( 'X', 'r', 'S', 'X', 'S', '-', 'X' ),
	( 'X', 'f', 'S', 'X', 'S', '-', 'X' ),
	( 'X', 'X', 'S', 'r', 'S', '-', 'X' ),
	( 'X', 'X', 'S', 'f', 'S', '-', 'X' ),
	( 'X', 'X', 'S', 'X', 'S', '-', 'S' ),
	( 'S', 'S', 'r', 'X', 'S', '-', 'X' ),
	( 'S', 'S', 'f', 'X', 'S', '-', 'X' ),
	( 'S', 'S', 'X', 'r', 'S', '-', 'X' ),
	( 'S', 'S', 'X', 'f', 'S', '-', 'X' ),
	( 'S', 'S', 'X', 'X', 'S', '-', 'S' ),
	( 'r', 'S', 'X', 'X', 'S', '-', 'X' ),
	( 'f', 'S', 'X', 'X', 'S', '-', 'X' ),
	( 'X', 'S', 'r', 'X', 'S', '-', 'X' ),
	( 'X', 'S', 'f', 'X', 'S', '-', 'X' ),
	( 'X', 'S', 'X', 'r', 'S', '-', 'X' ),
	( 'X', 'S', 'X', 'f', 'S', '-', 'X' ),
	( 'X', 'S', 'X', 'X', 'S', '-', 'S' ),
	( 'S', 'r', 'X', 'X', 'S', '-', 'X' ),
	( 'S', 'f', 'X', 'X', 'S', '-', 'X' ),
	( 'S', 'X', 'r', 'X', 'S', '-', 'X' ),
	( 'S', 'X', 'f', 'X', 'S', '-', 'X' ),
	( 'S', 'X', 'X', 'r', 'S', '-', 'X' ),
	( 'S', 'X', 'X', 'f', 'S', '-', 'X' ),
	( 'S', 'X', 'X', 'X', 'S', '-', 'S' ),
	( 'r', 'X', 'X', 'X', 'S', '-', 'X' ),
	( 'f', 'X', 'X', 'X', 'S', '-', 'X' ),
	( 'X', 'r', 'X', 'X', 'S', '-', 'X' ),
	( 'X', 'f', 'X', 'X', 'S', '-', 'X' ),
	( 'X', 'X', 'r', 'X', 'S', '-', 'X' ),
	( 'X', 'X', 'f', 'X', 'S', '-', 'X' ),
	( 'X', 'X', 'X', 'r', 'S', '-', 'X' ),
	( 'X', 'X', 'X', 'f', 'S', '-', 'X' ),
	( 'X', 'X', 'X', 'X', 'S', '-', 'S' ),
	( 'S', 'S', 'S', 'S', 'r', '-', 'X' ),
	( 'S', 'S', 'S', 'S', 'f', '-', 'X' ),
	( 'S', 'S', 'S', 'S', 'X', '-', 'S' ),
	( 'r', 'S', 'S', 'S', 'X', '-', 'X' ),
	( 'f', 'S', 'S', 'S', 'X', '-', 'X' ),
	( 'X', 'S', 'S', 'S', 'r', '-', 'X' ),
	( 'X', 'S', 'S', 'S', 'f', '-', 'X' ),
	( 'X', 'S', 'S', 'S', 'X', '-', 'S' ),
	( 'S', 'r', 'S', 'S', 'X', '-', 'X' ),
	( 'S', 'f', 'S', 'S', 'X', '-', 'X' ),
	( 'S', 'X', 'S', 'S', 'r', '-', 'X' ),
	( 'S', 'X', 'S', 'S', 'f', '-', 'X' ),
	( 'S', 'X', 'S', 'S', 'X', '-', 'S' ),
	( 'r', 'X', 'S', 'S', 'X', '-', 'X' ),
	( 'f', 'X', 'S', 'S', 'X', '-', 'X' ),
	( 'X', 'r', 'S', 'S', 'X', '-', 'X' ),
	( 'X', 'f', 'S', 'S', 'X', '-', 'X' ),
	( 'X', 'X', 'S', 'S', 'r', '-', 'X' ),
	( 'X', 'X', 'S', 'S', 'f', '-', 'X' ),
	( 'X', 'X', 'S', 'S', 'X', '-', 'S' ),
	( 'S', 'S', 'r', 'S', 'X', '-', 'X' ),
	( 'S', 'S', 'f', 'S', 'X', '-', 'X' ),
	( 'S', 'S', 'X', 'S', 'r', '-', 'X' ),
	( 'S', 'S', 'X', 'S', 'f', '-', 'X' ),
	( 'S', 'S', 'X', 'S', 'X', '-', 'S' ),
	( 'r', 'S', 'X', 'S', 'X', '-', 'X' ),
	( 'f', 'S', 'X', 'S', 'X', '-', 'X' ),
	( 'X', 'S', 'r', 'S', 'X', '-', 'X' ),
	( 'X', 'S', 'f', 'S', 'X', '-', 'X' ),
	( 'X', 'S', 'X', 'S', 'r', '-', 'X' ),
	( 'X', 'S', 'X', 'S', 'f', '-', 'X' ),
	( 'X', 'S', 'X', 'S', 'X', '-', 'S' ),
	( 'S', 'r', 'X', 'S', 'X', '-', 'X' ),
	( 'S', 'f', 'X', 'S', 'X', '-', 'X' ),
	( 'S', 'X', 'r', 'S', 'X', '-', 'X' ),
	( 'S', 'X', 'f', 'S', 'X', '-', 'X' ),
	( 'S', 'X', 'X', 'S', 'r', '-', 'X' ),
	( 'S', 'X', 'X', 'S', 'f', '-', 'X' ),
	( 'S', 'X', 'X', 'S', 'X', '-', 'S' ),
	( 'r', 'X', 'X', 'S', 'X', '-', 'X' ),
	( 'f', 'X', 'X', 'S', 'X', '-', 'X' ),
	( 'X', 'r', 'X', 'S', 'X', '-', 'X' ),
	( 'X', 'f', 'X', 'S', 'X', '-', 'X' ),
	( 'X', 'X', 'r', 'S', 'X', '-', 'X' ),
	( 'X', 'X', 'f', 'S', 'X', '-', 'X' ),
	( 'X', 'X', 'X', 'S', 'r', '-', 'X' ),
	( 'X', 'X', 'X', 'S', 'f', '-', 'X' ),
	( 'X', 'X', 'X', 'S', 'X', '-', 'S' ),
	( 'S', 'S', 'S', 'r', 'X', '-', 'X' ),
	( 'S', 'S', 'S', 'f', 'X', '-', 'X' ),
	( 'S', 'S', 'S', 'X', 'r', '-', 'X' ),
	( 'S', 'S', 'S', 'X', 'f', '-', 'X' ),
	( 'S', 'S', 'S', 'X', 'X', '-', 'S' ),
	( 'r', 'S', 'S', 'X', 'X', '-', 'X' ),
	( 'f', 'S', 'S', 'X', 'X', '-', 'X' ),
	( 'X', 'S', 'S', 'r', 'X', '-', 'X' ),
	( 'X', 'S', 'S', 'f', 'X', '-', 'X' ),
	( 'X', 'S', 'S', 'X', 'r', '-', 'X' ),
	( 'X', 'S', 'S', 'X', 'f', '-', 'X' ),
	( 'X', 'S', 'S', 'X', 'X', '-', 'S' ),
	( 'S', 'r', 'S', 'X', 'X', '-', 'X' ),
	( 'S', 'f', 'S', 'X', 'X', '-', 'X' ),
	( 'S', 'X', 'S', 'r', 'X', '-', 'X' ),
	( 'S', 'X', 'S', 'f', 'X', '-', 'X' ),
	( 'S', 'X', 'S', 'X', 'r', '-', 'X' ),
	( 'S', 'X', 'S', 'X', 'f', '-', 'X' ),
	( 'S', 'X', 'S', 'X', 'X', '-', 'S' ),
	( 'r', 'X', 'S', 'X', 'X', '-', 'X' ),
	( 'f', 'X', 'S', 'X', 'X', '-', 'X' ),
	( 'X', 'r', 'S', 'X', 'X', '-', 'X' ),
	( 'X', 'f', 'S', 'X', 'X', '-', 'X' ),
	( 'X', 'X', 'S', 'r', 'X', '-', 'X' ),
	( 'X', 'X', 'S', 'f', 'X', '-', 'X' ),
	( 'X', 'X', 'S', 'X', 'r', '-', 'X' ),
	( 'X', 'X', 'S', 'X', 'f', '-', 'X' ),
	( 'X', 'X', 'S', 'X', 'X', '-', 'S' ),
	( 'S', 'S', 'r', 'X', 'X', '-', 'X' ),
	( 'S', 'S', 'f', 'X', 'X', '-', 'X' ),
	( 'S', 'S', 'X', 'r', 'X', '-', 'X' ),
	( 'S', 'S', 'X', 'f', 'X', '-', 'X' ),
	( 'S', 'S', 'X', 'X', 'r', '-', 'X' ),
	( 'S', 'S', 'X', 'X', 'f', '-', 'X' ),
	( 'S', 'S', 'X', 'X', 'X', '-', 'S' ),
	( 'r', 'S', 'X', 'X', 'X', '-', 'X' ),
	( 'f', 'S', 'X', 'X', 'X', '-', 'X' ),
	( 'X', 'S', 'r', 'X', 'X', '-', 'X' ),
	( 'X', 'S', 'f', 'X', 'X', '-', 'X' ),
	( 'X', 'S', 'X', 'r', 'X', '-', 'X' ),
	( 'X', 'S', 'X', 'f', 'X', '-', 'X' ),
	( 'X', 'S', 'X', 'X', 'r', '-', 'X' ),
	( 'X', 'S', 'X', 'X', 'f', '-', 'X' ),
	( 'X', 'S', 'X', 'X', 'X', '-', 'S' ),
	( 'S', 'r', 'X', 'X', 'X', '-', 'X' ),
	( 'S', 'f', 'X', 'X', 'X', '-', 'X' ),
	( 'S', 'X', 'r', 'X', 'X', '-', 'X' ),
	( 'S', 'X', 'f', 'X', 'X', '-', 'X' ),
	( 'S', 'X', 'X', 'r', 'X', '-', 'X' ),
	( 'S', 'X', 'X', 'f', 'X', '-', 'X' ),
	( 'S', 'X', 'X', 'X', 'r', '-', 'X' ),
	( 'S', 'X', 'X', 'X', 'f', '-', 'X' ),
	( 'S', 'X', 'X', 'X', 'X', '-', 'S' ),
	( 'r', 'X', 'X', 'X', 'X', '-', 'X' ),
	( 'f', 'X', 'X', 'X', 'X', '-', 'X' ),
	( 'X', 'r', 'X', 'X', 'X', '-', 'X' ),
	( 'X', 'f', 'X', 'X', 'X', '-', 'X' ),
	( 'X', 'X', 'r', 'X', 'X', '-', 'X' ),
	( 'X', 'X', 'f', 'X', 'X', '-', 'X' ),
	( 'X', 'X', 'X', 'r', 'X', '-', 'X' ),
	( 'X', 'X', 'X', 'f', 'X', '-', 'X' ),
	( 'X', 'X', 'X', 'X', 'r', '-', 'X' ),
	( 'X', 'X', 'X', 'X', 'f', '-', 'X' ),
	( 'X', 'X', 'X', 'X', 'X', '-', 'S' ) );


	-------------------------------------------------------------------------------
	--State Table Declaration
	-------------------------------------------------------------------------------
	CONSTANT rsfftab : VitalStateTableType := (
	-- CLK RE SE S R lstSt Q
	( '-', '-', '-', '0', '1', '-', '1' ),
	( '-', '-', '-', '1', '0', '-', '0' ),
	( '-', '1', '1', '/', '1', '-', 'S' ),
	( '-', '1', '1', '^', '1', '-', 'S' ),
	( '-', '1', '1', '1', '/', '-', 'S' ),
	( '-', '1', '1', '1', '^', '-', 'S' ),
	( '/', '0', '0', '1', '1', '-', 'S' ),
	( '/', '0', '1', '1', '1', '-', '1' ),
	( '/', '1', '0', '1', '1', '-', '0' ),
	( '\', '-', '-', '-', '-', '-', 'S' ),
	( 'R', '0', '0', '1', '1', '-', 'S' ),
	( 'R', '0', '-', '1', '-', '0', 'S' ),
	( 'R', '-', '0', '-', '1', '1', 'S' ),
	( 'v', '-', '-', '-', '-', '-', 'S' ),
	( 'f', '0', '0', '1', '1', '-', 'S' ),
	( 'f', '0', '-', '1', '-', '0', 'S' ),
	( 'f', '-', '0', '-', '1', '1', 'S' ),
	( 'X', '*', '0', '-', '1', '1', 'S' ),
	( 'X', '0', '*', '1', '-', '0', 'S' ),
	( 'S', 'S', 'S', 'S', 'S', '-', 'S' ),
	( 'r', 'S', 'S', 'S', 'S', '-', 'X' ),
	( 'f', 'S', 'S', 'S', 'S', '-', 'X' ),
	( 'X', 'S', 'S', 'S', 'S', '-', 'S' ),
	( 'S', 'r', 'S', 'S', 'S', '-', 'X' ),
	( 'S', 'f', 'S', 'S', 'S', '-', 'X' ),
	( 'S', 'X', 'S', 'S', 'S', '-', 'S' ),
	( 'r', 'X', 'S', 'S', 'S', '-', 'X' ),
	( 'f', 'X', 'S', 'S', 'S', '-', 'X' ),
	( 'X', 'r', 'S', 'S', 'S', '-', 'X' ),
	( 'X', 'f', 'S', 'S', 'S', '-', 'X' ),
	( 'X', 'X', 'S', 'S', 'S', '-', 'S' ),
	( 'S', 'S', 'r', 'S', 'S', '-', 'X' ),
	( 'S', 'S', 'f', 'S', 'S', '-', 'X' ),
	( 'S', 'S', 'X', 'S', 'S', '-', 'S' ),
	( 'r', 'S', 'X', 'S', 'S', '-', 'X' ),
	( 'f', 'S', 'X', 'S', 'S', '-', 'X' ),
	( 'X', 'S', 'r', 'S', 'S', '-', 'X' ),
	( 'X', 'S', 'f', 'S', 'S', '-', 'X' ),
	( 'X', 'S', 'X', 'S', 'S', '-', 'S' ),
	( 'S', 'r', 'X', 'S', 'S', '-', 'X' ),
	( 'S', 'f', 'X', 'S', 'S', '-', 'X' ),
	( 'S', 'X', 'r', 'S', 'S', '-', 'X' ),
	( 'S', 'X', 'f', 'S', 'S', '-', 'X' ),
	( 'S', 'X', 'X', 'S', 'S', '-', 'S' ),
	( 'r', 'X', 'X', 'S', 'S', '-', 'X' ),
	( 'f', 'X', 'X', 'S', 'S', '-', 'X' ),
	( 'X', 'r', 'X', 'S', 'S', '-', 'X' ),
	( 'X', 'f', 'X', 'S', 'S', '-', 'X' ),
	( 'X', 'X', 'r', 'S', 'S', '-', 'X' ),
	( 'X', 'X', 'f', 'S', 'S', '-', 'X' ),
	( 'X', 'X', 'X', 'S', 'S', '-', 'S' ),
	( 'S', 'S', 'S', 'r', 'S', '-', 'X' ),
	( 'S', 'S', 'S', 'f', 'S', '-', 'X' ),
	( 'S', 'S', 'S', 'X', 'S', '-', 'S' ),
	( 'r', 'S', 'S', 'X', 'S', '-', 'X' ),
	( 'f', 'S', 'S', 'X', 'S', '-', 'X' ),
	( 'X', 'S', 'S', 'r', 'S', '-', 'X' ),
	( 'X', 'S', 'S', 'f', 'S', '-', 'X' ),
	( 'X', 'S', 'S', 'X', 'S', '-', 'S' ),
	( 'S', 'r', 'S', 'X', 'S', '-', 'X' ),
	( 'S', 'f', 'S', 'X', 'S', '-', 'X' ),
	( 'S', 'X', 'S', 'r', 'S', '-', 'X' ),
	( 'S', 'X', 'S', 'f', 'S', '-', 'X' ),
	( 'S', 'X', 'S', 'X', 'S', '-', 'S' ),
	( 'r', 'X', 'S', 'X', 'S', '-', 'X' ),
	( 'f', 'X', 'S', 'X', 'S', '-', 'X' ),
	( 'X', 'r', 'S', 'X', 'S', '-', 'X' ),
	( 'X', 'f', 'S', 'X', 'S', '-', 'X' ),
	( 'X', 'X', 'S', 'r', 'S', '-', 'X' ),
	( 'X', 'X', 'S', 'f', 'S', '-', 'X' ),
	( 'X', 'X', 'S', 'X', 'S', '-', 'S' ),
	( 'S', 'S', 'r', 'X', 'S', '-', 'X' ),
	( 'S', 'S', 'f', 'X', 'S', '-', 'X' ),
	( 'S', 'S', 'X', 'r', 'S', '-', 'X' ),
	( 'S', 'S', 'X', 'f', 'S', '-', 'X' ),
	( 'S', 'S', 'X', 'X', 'S', '-', 'S' ),
	( 'r', 'S', 'X', 'X', 'S', '-', 'X' ),
	( 'f', 'S', 'X', 'X', 'S', '-', 'X' ),
	( 'X', 'S', 'r', 'X', 'S', '-', 'X' ),
	( 'X', 'S', 'f', 'X', 'S', '-', 'X' ),
	( 'X', 'S', 'X', 'r', 'S', '-', 'X' ),
	( 'X', 'S', 'X', 'f', 'S', '-', 'X' ),
	( 'X', 'S', 'X', 'X', 'S', '-', 'S' ),
	( 'S', 'r', 'X', 'X', 'S', '-', 'X' ),
	( 'S', 'f', 'X', 'X', 'S', '-', 'X' ),
	( 'S', 'X', 'r', 'X', 'S', '-', 'X' ),
	( 'S', 'X', 'f', 'X', 'S', '-', 'X' ),
	( 'S', 'X', 'X', 'r', 'S', '-', 'X' ),
	( 'S', 'X', 'X', 'f', 'S', '-', 'X' ),
	( 'S', 'X', 'X', 'X', 'S', '-', 'S' ),
	( 'r', 'X', 'X', 'X', 'S', '-', 'X' ),
	( 'f', 'X', 'X', 'X', 'S', '-', 'X' ),
	( 'X', 'r', 'X', 'X', 'S', '-', 'X' ),
	( 'X', 'f', 'X', 'X', 'S', '-', 'X' ),
	( 'X', 'X', 'r', 'X', 'S', '-', 'X' ),
	( 'X', 'X', 'f', 'X', 'S', '-', 'X' ),
	( 'X', 'X', 'X', 'r', 'S', '-', 'X' ),
	( 'X', 'X', 'X', 'f', 'S', '-', 'X' ),
	( 'X', 'X', 'X', 'X', 'S', '-', 'S' ),
	( 'S', 'S', 'S', 'S', '/', '-', 'S' ),----
	( 'S', 'S', 'S', '/', 'S', '-', 'S' ),----
	( 'S', 'S', 'S', 'S', 'r', '-', 'X' ),----
	( 'S', 'S', 'S', 'S', 'f', '-', 'X' ),
	( 'S', 'S', 'S', 'S', 'X', '-', 'S' ),
	( 'r', 'S', 'S', 'S', 'X', '-', 'X' ),
	( 'f', 'S', 'S', 'S', 'X', '-', 'X' ),
	( 'X', 'S', 'S', 'S', 'r', '-', 'X' ),
	( 'X', 'S', 'S', 'S', 'f', '-', 'X' ),
	( 'X', 'S', 'S', 'S', 'X', '-', 'S' ),
	( 'S', 'r', 'S', 'S', 'X', '-', 'X' ),
	( 'S', 'f', 'S', 'S', 'X', '-', 'X' ),
	( 'S', 'X', 'S', 'S', 'r', '-', 'X' ),
	( 'S', 'X', 'S', 'S', 'f', '-', 'X' ),
	( 'S', 'X', 'S', 'S', 'X', '-', 'S' ),
	( 'r', 'X', 'S', 'S', 'X', '-', 'X' ),
	( 'f', 'X', 'S', 'S', 'X', '-', 'X' ),
	( 'X', 'r', 'S', 'S', 'X', '-', 'X' ),
	( 'X', 'f', 'S', 'S', 'X', '-', 'X' ),
	( 'X', 'X', 'S', 'S', 'r', '-', 'X' ),
	( 'X', 'X', 'S', 'S', 'f', '-', 'X' ),
	( 'X', 'X', 'S', 'S', 'X', '-', 'S' ),
	( 'S', 'S', 'r', 'S', 'X', '-', 'X' ),
	( 'S', 'S', 'f', 'S', 'X', '-', 'X' ),
	( 'S', 'S', 'X', 'S', 'r', '-', 'X' ),
	( 'S', 'S', 'X', 'S', 'f', '-', 'X' ),
	( 'S', 'S', 'X', 'S', 'X', '-', 'S' ),
	( 'r', 'S', 'X', 'S', 'X', '-', 'X' ),
	( 'f', 'S', 'X', 'S', 'X', '-', 'X' ),
	( 'X', 'S', 'r', 'S', 'X', '-', 'X' ),
	( 'X', 'S', 'f', 'S', 'X', '-', 'X' ),
	( 'X', 'S', 'X', 'S', 'r', '-', 'X' ),
	( 'X', 'S', 'X', 'S', 'f', '-', 'X' ),
	( 'X', 'S', 'X', 'S', 'X', '-', 'S' ),
	( 'S', 'r', 'X', 'S', 'X', '-', 'X' ),
	( 'S', 'f', 'X', 'S', 'X', '-', 'X' ),
	( 'S', 'X', 'r', 'S', 'X', '-', 'X' ),
	( 'S', 'X', 'f', 'S', 'X', '-', 'X' ),
	( 'S', 'X', 'X', 'S', 'r', '-', 'X' ),
	( 'S', 'X', 'X', 'S', 'f', '-', 'X' ),
	( 'S', 'X', 'X', 'S', 'X', '-', 'S' ),
	( 'r', 'X', 'X', 'S', 'X', '-', 'X' ),
	( 'f', 'X', 'X', 'S', 'X', '-', 'X' ),
	( 'X', 'r', 'X', 'S', 'X', '-', 'X' ),
	( 'X', 'f', 'X', 'S', 'X', '-', 'X' ),
	( 'X', 'X', 'r', 'S', 'X', '-', 'X' ),
	( 'X', 'X', 'f', 'S', 'X', '-', 'X' ),
	( 'X', 'X', 'X', 'S', 'r', '-', 'X' ),
	( 'X', 'X', 'X', 'S', 'f', '-', 'X' ),
	( 'X', 'X', 'X', 'S', 'X', '-', 'S' ),
	( 'S', 'S', 'S', 'r', 'X', '-', 'X' ),
	( 'S', 'S', 'S', 'f', 'X', '-', 'X' ),
	( 'S', 'S', 'S', 'X', 'r', '-', 'X' ),
	( 'S', 'S', 'S', 'X', 'f', '-', 'X' ),
	( 'S', 'S', 'S', 'X', 'X', '-', 'S' ),
	( 'r', 'S', 'S', 'X', 'X', '-', 'X' ),
	( 'f', 'S', 'S', 'X', 'X', '-', 'X' ),
	( 'X', 'S', 'S', 'r', 'X', '-', 'X' ),
	( 'X', 'S', 'S', 'f', 'X', '-', 'X' ),
	( 'X', 'S', 'S', 'X', 'r', '-', 'X' ),
	( 'X', 'S', 'S', 'X', 'f', '-', 'X' ),
	( 'X', 'S', 'S', 'X', 'X', '-', 'S' ),
	( 'S', 'r', 'S', 'X', 'X', '-', 'X' ),
	( 'S', 'f', 'S', 'X', 'X', '-', 'X' ),
	( 'S', 'X', 'S', 'r', 'X', '-', 'X' ),
	( 'S', 'X', 'S', 'f', 'X', '-', 'X' ),
	( 'S', 'X', 'S', 'X', 'r', '-', 'X' ),
	( 'S', 'X', 'S', 'X', 'f', '-', 'X' ),
	( 'S', 'X', 'S', 'X', 'X', '-', 'S' ),
	( 'r', 'X', 'S', 'X', 'X', '-', 'X' ),
	( 'f', 'X', 'S', 'X', 'X', '-', 'X' ),
	( 'X', 'r', 'S', 'X', 'X', '-', 'X' ),
	( 'X', 'f', 'S', 'X', 'X', '-', 'X' ),
	( 'X', 'X', 'S', 'r', 'X', '-', 'X' ),
	( 'X', 'X', 'S', 'f', 'X', '-', 'X' ),
	( 'X', 'X', 'S', 'X', 'r', '-', 'X' ),
	( 'X', 'X', 'S', 'X', 'f', '-', 'X' ),
	( 'X', 'X', 'S', 'X', 'X', '-', 'S' ),
	( 'S', 'S', 'r', 'X', 'X', '-', 'X' ),
	( 'S', 'S', 'f', 'X', 'X', '-', 'X' ),
	( 'S', 'S', 'X', 'r', 'X', '-', 'X' ),
	( 'S', 'S', 'X', 'f', 'X', '-', 'X' ),
	( 'S', 'S', 'X', 'X', 'r', '-', 'X' ),
	( 'S', 'S', 'X', 'X', 'f', '-', 'X' ),
	( 'S', 'S', 'X', 'X', 'X', '-', 'S' ),
	( 'r', 'S', 'X', 'X', 'X', '-', 'X' ),
	( 'f', 'S', 'X', 'X', 'X', '-', 'X' ),
	( 'X', 'S', 'r', 'X', 'X', '-', 'X' ),
	( 'X', 'S', 'f', 'X', 'X', '-', 'X' ),
	( 'X', 'S', 'X', 'r', 'X', '-', 'X' ),
	( 'X', 'S', 'X', 'f', 'X', '-', 'X' ),
	( 'X', 'S', 'X', 'X', 'r', '-', 'X' ),
	( 'X', 'S', 'X', 'X', 'f', '-', 'X' ),
	( 'X', 'S', 'X', 'X', 'X', '-', 'S' ),
	( 'S', 'r', 'X', 'X', 'X', '-', 'X' ),
	( 'S', 'f', 'X', 'X', 'X', '-', 'X' ),
	( 'S', 'X', 'r', 'X', 'X', '-', 'X' ),
	( 'S', 'X', 'f', 'X', 'X', '-', 'X' ),
	( 'S', 'X', 'X', 'r', 'X', '-', 'X' ),
	( 'S', 'X', 'X', 'f', 'X', '-', 'X' ),
	( 'S', 'X', 'X', 'X', 'r', '-', 'X' ),
	( 'S', 'X', 'X', 'X', 'f', '-', 'X' ),
	( 'S', 'X', 'X', 'X', 'X', '-', 'S' ),
	( 'r', 'X', 'X', 'X', 'X', '-', 'X' ),
	( 'f', 'X', 'X', 'X', 'X', '-', 'X' ),
	( 'X', 'r', 'X', 'X', 'X', '-', 'X' ),
	( 'X', 'f', 'X', 'X', 'X', '-', 'X' ),
	( 'X', 'X', 'r', 'X', 'X', '-', 'X' ),
	( 'X', 'X', 'f', 'X', 'X', '-', 'X' ),
	( 'X', 'X', 'X', 'r', 'X', '-', 'X' ),
	( 'X', 'X', 'X', 'f', 'X', '-', 'X' ),
	( 'X', 'X', 'X', 'X', 'r', '-', 'X' ),
	( 'X', 'X', 'X', 'X', 'f', '-', 'X' ),
	( 'X', 'X', 'X', 'X', 'X', '-', 'S' ),
	( '-', '*', '-', '1', '1', '-', 'S' ),
	( '-', '-', '*', '1', '1', '-', 'S' ));


	-------------------------------------------------------------------------------
	--State Table Declaration
	-------------------------------------------------------------------------------
	CONSTANT tfftab : VitalStateTableType := (
	-- CLK T S R lstSt Q
	( '-', '-', '0', '1', '-', '1' ),
	( '-', '-', '1', '0', '-', '0' ),
	( 'X', '0', '1', '-', '0', 'S' ),
	( '-', '-', '*', '1', '1', '1' ),
	( '-', '-', '1', '*', '0', '0' ),
	( '/', '0', '1', '1', '-', 'S' ),
	( '/', '1', '1', '1', '1', '0' ),
	( '/', '1', '1', '1', '0', '1' ),
	( '\', '-', '-', '-', '-', 'S' ),
	( 'B', '*', '-', '-', '-', 'S' ),
	( 'R', '0', '1', '1', '-', 'S' ),
	( 'R', '0', '1', '-', '0', 'S' ),
	( 'R', '0', '-', '1', '1', 'S' ),
	( 'v', '-', '-', '-', '-', 'S' ),
	( 'f', '0', '1', '1', '-', 'S' ),
	( 'f', '-', '-', '1', '1', 'S' ),
	( 'S', 'S', 'S', 'S', '-', 'S' ),
	( 'r', 'S', 'S', 'S', '-', 'X' ),
	( 'f', 'S', 'S', 'S', '-', 'X' ),
	( 'X', 'S', 'S', 'S', '-', 'S' ),
	( 'S', 'r', 'S', 'S', '-', 'X' ),
	( 'S', 'f', 'S', 'S', '-', 'X' ),
	( 'S', 'X', 'S', 'S', '-', 'S' ),
	( 'r', 'X', 'S', 'S', '-', 'X' ),
	( 'f', 'X', 'S', 'S', '-', 'X' ),
	( 'X', 'r', 'S', 'S', '-', 'X' ),
	( 'X', 'f', 'S', 'S', '-', 'X' ),
	( 'X', 'X', 'S', 'S', '-', 'S' ),
	( 'S', 'S', 'r', 'S', '-', 'X' ),
	( 'S', 'S', 'f', 'S', '-', 'X' ),
	( 'S', 'S', 'X', 'S', '-', 'S' ),
	( 'r', 'S', 'X', 'S', '-', 'X' ),
	( 'f', 'S', 'X', 'S', '-', 'X' ),
	( 'X', 'S', 'r', 'S', '-', 'X' ),
	( 'X', 'S', 'f', 'S', '-', 'X' ),
	( 'X', 'S', 'X', 'S', '-', 'S' ),
	( 'S', 'r', 'X', 'S', '-', 'X' ),
	( 'S', 'f', 'X', 'S', '-', 'X' ),
	( 'S', 'X', 'r', 'S', '-', 'X' ),
	( 'S', 'X', 'f', 'S', '-', 'X' ),
	( 'S', 'X', 'X', 'S', '-', 'S' ),
	( 'r', 'X', 'X', 'S', '-', 'X' ),
	( 'f', 'X', 'X', 'S', '-', 'X' ),
	( 'X', 'r', 'X', 'S', '-', 'X' ),
	( 'X', 'f', 'X', 'S', '-', 'X' ),
	( 'X', 'X', 'r', 'S', '-', 'X' ),
	( 'X', 'X', 'f', 'S', '-', 'X' ),
	( 'X', 'X', 'X', 'S', '-', 'S' ),
	( 'S', 'S', 'S', 'r', '-', 'X' ),
	( 'S', 'S', 'S', 'f', '-', 'X' ),
	( 'S', 'S', 'S', 'X', '-', 'S' ),
	( 'r', 'S', 'S', 'X', '-', 'X' ),
	( 'f', 'S', 'S', 'X', '-', 'X' ),
	( 'X', 'S', 'S', 'r', '-', 'X' ),
	( 'X', 'S', 'S', 'f', '-', 'X' ),
	( 'X', 'S', 'S', 'X', '-', 'S' ),
	( 'S', 'r', 'S', 'X', '-', 'X' ),
	( 'S', 'f', 'S', 'X', '-', 'X' ),
	( 'S', 'X', 'S', 'r', '-', 'X' ),
	( 'S', 'X', 'S', 'f', '-', 'X' ),
	( 'S', 'X', 'S', 'X', '-', 'S' ),
	( 'r', 'X', 'S', 'X', '-', 'X' ),
	( 'f', 'X', 'S', 'X', '-', 'X' ),
	( 'X', 'r', 'S', 'X', '-', 'X' ),
	( 'X', 'f', 'S', 'X', '-', 'X' ),
	( 'X', 'X', 'S', 'r', '-', 'X' ),
	( 'X', 'X', 'S', 'f', '-', 'X' ),
	( 'X', 'X', 'S', 'X', '-', 'S' ),
	( 'S', 'S', 'r', 'X', '-', 'X' ),
	( 'S', 'S', 'f', 'X', '-', 'X' ),
	( 'S', 'S', 'X', 'r', '-', 'X' ),
	( 'S', 'S', 'X', 'f', '-', 'X' ),
	( 'S', 'S', 'X', 'X', '-', 'S' ),
	( 'r', 'S', 'X', 'X', '-', 'X' ),
	( 'f', 'S', 'X', 'X', '-', 'X' ),
	( 'X', 'S', 'r', 'X', '-', 'X' ),
	( 'X', 'S', 'f', 'X', '-', 'X' ),
	( 'X', 'S', 'X', 'r', '-', 'X' ),
	( 'X', 'S', 'X', 'f', '-', 'X' ),
	( 'X', 'S', 'X', 'X', '-', 'S' ),
	( 'S', 'r', 'X', 'X', '-', 'X' ),
	( 'S', 'f', 'X', 'X', '-', 'X' ),
	( 'S', 'X', 'r', 'X', '-', 'X' ),
	( 'S', 'X', 'f', 'X', '-', 'X' ),
	( 'S', 'X', 'X', 'r', '-', 'X' ),
	( 'S', 'X', 'X', 'f', '-', 'X' ),
	( 'S', 'X', 'X', 'X', '-', 'S' ),
	( 'r', 'X', 'X', 'X', '-', 'X' ),
	( 'f', 'X', 'X', 'X', '-', 'X' ),
	( 'X', 'r', 'X', 'X', '-', 'X' ),
	( 'X', 'f', 'X', 'X', '-', 'X' ),
	( 'X', 'X', 'r', 'X', '-', 'X' ),
	( 'X', 'X', 'f', 'X', '-', 'X' ),
	( 'X', 'X', 'X', 'r', '-', 'X' ),
	( 'X', 'X', 'X', 'f', '-', 'X' ),
	( 'X', 'X', 'X', 'X', '-', 'S' ) );


	-------------------------------------------------------------------------------
	--State Table Declaration
	-------------------------------------------------------------------------------
	CONSTANT dffcetab : VitalStateTableType := (
	-- D CLK R S CE lstSt Q
	( '-', '-', '0', '1', '-', '-', '0' ),
	( '-', '-', '1', '0', '-', '-', '1' ),
	( '-', '-', '1', '1', '0', '-', 'S' ),
	( '1', '/', '1', '-', '1', '-', '1' ),
	( '0', '/', '-', '1', '1', '-', '0' ),
	( '1', '-', '1', '*', '1', '1', '1' ),
	( '-', '0', '1', '*', '1', '1', '1' ),
	( '-', '1', '1', '*', '1', '1', '1' ),
	( '0', '-', '*', '1', '1', '0', '0' ),
	( '-', '0', '*', '1', '1', '0', '0' ),
	( '-', '1', '*', '1', '1', '0', '0' ),
	( '1', 'R', '1', '1', '1', '1', '1' ),
	( '0', 'R', '1', '1', '1', '0', '0' ),
	( '-', '\', '-', '-', '1', '-', 'S' ),
	( '-', 'v', '-', '-', '1', '-', 'S' ),
	( '0', 'r', '-', '-', '1', '0', 'S' ),
	( '0', 'f', '-', '-', '1', '0', 'S' ),
	( '1', 'r', '-', '-', '1', '1', 'S' ),
	( '1', 'f', '-', '-', '1', '1', 'S' ),
	( '*', '1', '-', '-', '1', '-', 'S' ),
	( '*', '0', '-', '-', '1', '-', 'S' ),
	( 'S', 'S', 'S', 'S', 'S', '-', 'S' ),
	( 'r', 'S', 'S', 'S', 'S', '-', 'X' ),
	( 'f', 'S', 'S', 'S', 'S', '-', 'X' ),
	( 'X', 'S', 'S', 'S', 'S', '-', 'S' ),
	( 'S', 'r', 'S', 'S', 'S', '-', 'X' ),
	( 'S', 'f', 'S', 'S', 'S', '-', 'X' ),
	( 'S', 'X', 'S', 'S', 'S', '-', 'S' ),
	( 'r', 'X', 'S', 'S', 'S', '-', 'X' ),
	( 'f', 'X', 'S', 'S', 'S', '-', 'X' ),
	( 'X', 'r', 'S', 'S', 'S', '-', 'X' ),
	( 'X', 'f', 'S', 'S', 'S', '-', 'X' ),
	( 'X', 'X', 'S', 'S', 'S', '-', 'S' ),
	( 'S', 'S', 'r', 'S', 'S', '-', 'X' ),
	( 'S', 'S', 'f', 'S', 'S', '-', 'X' ),
	( 'S', 'S', 'X', 'S', 'S', '-', 'S' ),
	( 'r', 'S', 'X', 'S', 'S', '-', 'X' ),
	( 'f', 'S', 'X', 'S', 'S', '-', 'X' ),
	( 'X', 'S', 'r', 'S', 'S', '-', 'X' ),
	( 'X', 'S', 'f', 'S', 'S', '-', 'X' ),
	( 'X', 'S', 'X', 'S', 'S', '-', 'S' ),
	( 'S', 'r', 'X', 'S', 'S', '-', 'X' ),
	( 'S', 'f', 'X', 'S', 'S', '-', 'X' ),
	( 'S', 'X', 'r', 'S', 'S', '-', 'X' ),
	( 'S', 'X', 'f', 'S', 'S', '-', 'X' ),
	( 'S', 'X', 'X', 'S', 'S', '-', 'S' ),
	( 'r', 'X', 'X', 'S', 'S', '-', 'X' ),
	( 'f', 'X', 'X', 'S', 'S', '-', 'X' ),
	( 'X', 'r', 'X', 'S', 'S', '-', 'X' ),
	( 'X', 'f', 'X', 'S', 'S', '-', 'X' ),
	( 'X', 'X', 'r', 'S', 'S', '-', 'X' ),
	( 'X', 'X', 'f', 'S', 'S', '-', 'X' ),
	( 'X', 'X', 'X', 'S', 'S', '-', 'S' ),
	( 'S', 'S', 'S', 'r', 'S', '-', 'X' ),
	( 'S', 'S', 'S', 'f', 'S', '-', 'X' ),
	( 'S', 'S', 'S', 'X', 'S', '-', 'S' ),
	( 'r', 'S', 'S', 'X', 'S', '-', 'X' ),
	( 'f', 'S', 'S', 'X', 'S', '-', 'X' ),
	( 'X', 'S', 'S', 'r', 'S', '-', 'X' ),
	( 'X', 'S', 'S', 'f', 'S', '-', 'X' ),
	( 'X', 'S', 'S', 'X', 'S', '-', 'S' ),
	( 'S', 'r', 'S', 'X', 'S', '-', 'X' ),
	( 'S', 'f', 'S', 'X', 'S', '-', 'X' ),
	( 'S', 'X', 'S', 'r', 'S', '-', 'X' ),
	( 'S', 'X', 'S', 'f', 'S', '-', 'X' ),
	( 'S', 'X', 'S', 'X', 'S', '-', 'S' ),
	( 'r', 'X', 'S', 'X', 'S', '-', 'X' ),
	( 'f', 'X', 'S', 'X', 'S', '-', 'X' ),
	( 'X', 'r', 'S', 'X', 'S', '-', 'X' ),
	( 'X', 'f', 'S', 'X', 'S', '-', 'X' ),
	( 'X', 'X', 'S', 'r', 'S', '-', 'X' ),
	( 'X', 'X', 'S', 'f', 'S', '-', 'X' ),
	( 'X', 'X', 'S', 'X', 'S', '-', 'S' ),
	( 'S', 'S', 'r', 'X', 'S', '-', 'X' ),
	( 'S', 'S', 'f', 'X', 'S', '-', 'X' ),
	( 'S', 'S', 'X', 'r', 'S', '-', 'X' ),
	( 'S', 'S', 'X', 'f', 'S', '-', 'X' ),
	( 'S', 'S', 'X', 'X', 'S', '-', 'S' ),
	( 'r', 'S', 'X', 'X', 'S', '-', 'X' ),
	( 'f', 'S', 'X', 'X', 'S', '-', 'X' ),
	( 'X', 'S', 'r', 'X', 'S', '-', 'X' ),
	( 'X', 'S', 'f', 'X', 'S', '-', 'X' ),
	( 'X', 'S', 'X', 'r', 'S', '-', 'X' ),
	( 'X', 'S', 'X', 'f', 'S', '-', 'X' ),
	( 'X', 'S', 'X', 'X', 'S', '-', 'S' ),
	( 'S', 'r', 'X', 'X', 'S', '-', 'X' ),
	( 'S', 'f', 'X', 'X', 'S', '-', 'X' ),
	( 'S', 'X', 'r', 'X', 'S', '-', 'X' ),
	( 'S', 'X', 'f', 'X', 'S', '-', 'X' ),
	( 'S', 'X', 'X', 'r', 'S', '-', 'X' ),
	( 'S', 'X', 'X', 'f', 'S', '-', 'X' ),
	( 'S', 'X', 'X', 'X', 'S', '-', 'S' ),
	( 'r', 'X', 'X', 'X', 'S', '-', 'X' ),
	( 'f', 'X', 'X', 'X', 'S', '-', 'X' ),
	( 'X', 'r', 'X', 'X', 'S', '-', 'X' ),
	( 'X', 'f', 'X', 'X', 'S', '-', 'X' ),
	( 'X', 'X', 'r', 'X', 'S', '-', 'X' ),
	( 'X', 'X', 'f', 'X', 'S', '-', 'X' ),
	( 'X', 'X', 'X', 'r', 'S', '-', 'X' ),
	( 'X', 'X', 'X', 'f', 'S', '-', 'X' ),
	( 'X', 'X', 'X', 'X', 'S', '-', 'S' ),
	( 'S', 'S', 'S', 'S', 'r', '-', 'X' ),
	( 'S', 'S', 'S', 'S', 'f', '-', 'X' ),
	( 'S', 'S', 'S', 'S', 'X', '-', 'S' ),
	( 'r', 'S', 'S', 'S', 'X', '-', 'X' ),
	( 'f', 'S', 'S', 'S', 'X', '-', 'X' ),
	( 'X', 'S', 'S', 'S', 'r', '-', 'X' ),
	( 'X', 'S', 'S', 'S', 'f', '-', 'X' ),
	( 'X', 'S', 'S', 'S', 'X', '-', 'S' ),
	( 'S', 'r', 'S', 'S', 'X', '-', 'X' ),
	( 'S', 'f', 'S', 'S', 'X', '-', 'X' ),
	( 'S', 'X', 'S', 'S', 'r', '-', 'X' ),
	( 'S', 'X', 'S', 'S', 'f', '-', 'X' ),
	( 'S', 'X', 'S', 'S', 'X', '-', 'S' ),
	( 'r', 'X', 'S', 'S', 'X', '-', 'X' ),
	( 'f', 'X', 'S', 'S', 'X', '-', 'X' ),
	( 'X', 'r', 'S', 'S', 'X', '-', 'X' ),
	( 'X', 'f', 'S', 'S', 'X', '-', 'X' ),
	( 'X', 'X', 'S', 'S', 'r', '-', 'X' ),
	( 'X', 'X', 'S', 'S', 'f', '-', 'X' ),
	( 'X', 'X', 'S', 'S', 'X', '-', 'S' ),
	( 'S', 'S', 'r', 'S', 'X', '-', 'X' ),
	( 'S', 'S', 'f', 'S', 'X', '-', 'X' ),
	( 'S', 'S', 'X', 'S', 'r', '-', 'X' ),
	( 'S', 'S', 'X', 'S', 'f', '-', 'X' ),
	( 'S', 'S', 'X', 'S', 'X', '-', 'S' ),
	( 'r', 'S', 'X', 'S', 'X', '-', 'X' ),
	( 'f', 'S', 'X', 'S', 'X', '-', 'X' ),
	( 'X', 'S', 'r', 'S', 'X', '-', 'X' ),
	( 'X', 'S', 'f', 'S', 'X', '-', 'X' ),
	( 'X', 'S', 'X', 'S', 'r', '-', 'X' ),
	( 'X', 'S', 'X', 'S', 'f', '-', 'X' ),
	( 'X', 'S', 'X', 'S', 'X', '-', 'S' ),
	( 'S', 'r', 'X', 'S', 'X', '-', 'X' ),
	( 'S', 'f', 'X', 'S', 'X', '-', 'X' ),
	( 'S', 'X', 'r', 'S', 'X', '-', 'X' ),
	( 'S', 'X', 'f', 'S', 'X', '-', 'X' ),
	( 'S', 'X', 'X', 'S', 'r', '-', 'X' ),
	( 'S', 'X', 'X', 'S', 'f', '-', 'X' ),
	( 'S', 'X', 'X', 'S', 'X', '-', 'S' ),
	( 'r', 'X', 'X', 'S', 'X', '-', 'X' ),
	( 'f', 'X', 'X', 'S', 'X', '-', 'X' ),
	( 'X', 'r', 'X', 'S', 'X', '-', 'X' ),
	( 'X', 'f', 'X', 'S', 'X', '-', 'X' ),
	( 'X', 'X', 'r', 'S', 'X', '-', 'X' ),
	( 'X', 'X', 'f', 'S', 'X', '-', 'X' ),
	( 'X', 'X', 'X', 'S', 'r', '-', 'X' ),
	( 'X', 'X', 'X', 'S', 'f', '-', 'X' ),
	( 'X', 'X', 'X', 'S', 'X', '-', 'S' ),
	( 'S', 'S', 'S', 'r', 'X', '-', 'X' ),
	( 'S', 'S', 'S', 'f', 'X', '-', 'X' ),
	( 'S', 'S', 'S', 'X', 'r', '-', 'X' ),
	( 'S', 'S', 'S', 'X', 'f', '-', 'X' ),
	( 'S', 'S', 'S', 'X', 'X', '-', 'S' ),
	( 'r', 'S', 'S', 'X', 'X', '-', 'X' ),
	( 'f', 'S', 'S', 'X', 'X', '-', 'X' ),
	( 'X', 'S', 'S', 'r', 'X', '-', 'X' ),
	( 'X', 'S', 'S', 'f', 'X', '-', 'X' ),
	( 'X', 'S', 'S', 'X', 'r', '-', 'X' ),
	( 'X', 'S', 'S', 'X', 'f', '-', 'X' ),
	( 'X', 'S', 'S', 'X', 'X', '-', 'S' ),
	( 'S', 'r', 'S', 'X', 'X', '-', 'X' ),
	( 'S', 'f', 'S', 'X', 'X', '-', 'X' ),
	( 'S', 'X', 'S', 'r', 'X', '-', 'X' ),
	( 'S', 'X', 'S', 'f', 'X', '-', 'X' ),
	( 'S', 'X', 'S', 'X', 'r', '-', 'X' ),
	( 'S', 'X', 'S', 'X', 'f', '-', 'X' ),
	( 'S', 'X', 'S', 'X', 'X', '-', 'S' ),
	( 'r', 'X', 'S', 'X', 'X', '-', 'X' ),
	( 'f', 'X', 'S', 'X', 'X', '-', 'X' ),
	( 'X', 'r', 'S', 'X', 'X', '-', 'X' ),
	( 'X', 'f', 'S', 'X', 'X', '-', 'X' ),
	( 'X', 'X', 'S', 'r', 'X', '-', 'X' ),
	( 'X', 'X', 'S', 'f', 'X', '-', 'X' ),
	( 'X', 'X', 'S', 'X', 'r', '-', 'X' ),
	( 'X', 'X', 'S', 'X', 'f', '-', 'X' ),
	( 'X', 'X', 'S', 'X', 'X', '-', 'S' ),
	( 'S', 'S', 'r', 'X', 'X', '-', 'X' ),
	( 'S', 'S', 'f', 'X', 'X', '-', 'X' ),
	( 'S', 'S', 'X', 'r', 'X', '-', 'X' ),
	( 'S', 'S', 'X', 'f', 'X', '-', 'X' ),
	( 'S', 'S', 'X', 'X', 'r', '-', 'X' ),
	( 'S', 'S', 'X', 'X', 'f', '-', 'X' ),
	( 'S', 'S', 'X', 'X', 'X', '-', 'S' ),
	( 'r', 'S', 'X', 'X', 'X', '-', 'X' ),
	( 'f', 'S', 'X', 'X', 'X', '-', 'X' ),
	( 'X', 'S', 'r', 'X', 'X', '-', 'X' ),
	( 'X', 'S', 'f', 'X', 'X', '-', 'X' ),
	( 'X', 'S', 'X', 'r', 'X', '-', 'X' ),
	( 'X', 'S', 'X', 'f', 'X', '-', 'X' ),
	( 'X', 'S', 'X', 'X', 'r', '-', 'X' ),
	( 'X', 'S', 'X', 'X', 'f', '-', 'X' ),
	( 'X', 'S', 'X', 'X', 'X', '-', 'S' ),
	( 'S', 'r', 'X', 'X', 'X', '-', 'X' ),
	( 'S', 'f', 'X', 'X', 'X', '-', 'X' ),
	( 'S', 'X', 'r', 'X', 'X', '-', 'X' ),
	( 'S', 'X', 'f', 'X', 'X', '-', 'X' ),
	( 'S', 'X', 'X', 'r', 'X', '-', 'X' ),
	( 'S', 'X', 'X', 'f', 'X', '-', 'X' ),
	( 'S', 'X', 'X', 'X', 'r', '-', 'X' ),
	( 'S', 'X', 'X', 'X', 'f', '-', 'X' ),
	( 'S', 'X', 'X', 'X', 'X', '-', 'S' ),
	( 'r', 'X', 'X', 'X', 'X', '-', 'X' ),
	( 'f', 'X', 'X', 'X', 'X', '-', 'X' ),
	( 'X', 'r', 'X', 'X', 'X', '-', 'X' ),
	( 'X', 'f', 'X', 'X', 'X', '-', 'X' ),
	( 'X', 'X', 'r', 'X', 'X', '-', 'X' ),
	( 'X', 'X', 'f', 'X', 'X', '-', 'X' ),
	( 'X', 'X', 'X', 'r', 'X', '-', 'X' ),
	( 'X', 'X', 'X', 'f', 'X', '-', 'X' ),
	( 'X', 'X', 'X', 'X', 'r', '-', 'X' ),
	( 'X', 'X', 'X', 'X', 'f', '-', 'X' ),
	( '-', '-', '1', '1', '*', '-', 'S' ),
	( 'X', 'X', 'X', 'X', 'X', '-', 'S' ) );


end VLOGTOVITAL_TABLES;
----- VITAL model for cell AND10 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AND10 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_I0_O                       :	VitalDelayType01 := (3.050 ns, 3.050 ns);
      tpd_I1_O                       :	VitalDelayType01 := (3.050 ns, 3.050 ns);
      tpd_I2_O                       :	VitalDelayType01 := (3.050 ns, 3.050 ns);
      tpd_I3_O                       :	VitalDelayType01 := (3.050 ns, 3.050 ns);
      tpd_I4_O                       :	VitalDelayType01 := (3.050 ns, 3.050 ns);
      tpd_I5_O                       :	VitalDelayType01 := (3.050 ns, 3.050 ns);
      tpd_I6_O                       :	VitalDelayType01 := (3.050 ns, 3.050 ns);
      tpd_I7_O                       :	VitalDelayType01 := (3.050 ns, 3.050 ns);
      tpd_I8_O                       :	VitalDelayType01 := (3.050 ns, 3.050 ns);
      tpd_I9_O                       :	VitalDelayType01 := (3.050 ns, 3.050 ns);
      tipd_I0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I2                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I3                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I4                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I5                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I6                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I7                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I8                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I9                        :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      I0                             :	in    STD_ULOGIC;
      I1                             :	in    STD_ULOGIC;
      I2                             :	in    STD_ULOGIC;
      I3                             :	in    STD_ULOGIC;
      I4                             :	in    STD_ULOGIC;
      I5                             :	in    STD_ULOGIC;
      I6                             :	in    STD_ULOGIC;
      I7                             :	in    STD_ULOGIC;
      I8                             :	in    STD_ULOGIC;
      I9                             :	in    STD_ULOGIC;
      O                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AND10 : entity is TRUE;
end AND10;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
 
library VF1;
architecture VITAL_VF of AND10 is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL I0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I1_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I2_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I3_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I4_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I5_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I6_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I7_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I8_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I9_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (I0_ipd, I0, tipd_I0);
   VitalWireDelay (I1_ipd, I1, tipd_I1);
   VitalWireDelay (I2_ipd, I2, tipd_I2);
   VitalWireDelay (I3_ipd, I3, tipd_I3);
   VitalWireDelay (I4_ipd, I4, tipd_I4);
   VitalWireDelay (I5_ipd, I5, tipd_I5);
   VitalWireDelay (I6_ipd, I6, tipd_I6);
   VitalWireDelay (I7_ipd, I7, tipd_I7);
   VitalWireDelay (I8_ipd, I8, tipd_I8);
   VitalWireDelay (I9_ipd, I9, tipd_I9);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (I0_ipd, I1_ipd, I2_ipd, I3_ipd, I4_ipd, I5_ipd, I6_ipd, I7_ipd, I8_ipd, I9_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS O_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE O_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      O_zd :=
       (I1_ipd) AND (I0_ipd) AND (I2_ipd) AND (I3_ipd) AND (I4_ipd) AND
         (I5_ipd) AND (I6_ipd) AND (I7_ipd) AND (I8_ipd) AND (I9_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => O,
       GlitchData => O_GlitchData,
       OutSignalName => "O",
       OutTemp => O_zd,
       Paths => (0 => (I0_ipd'last_event, tpd_I0_O, TRUE),
                 1 => (I1_ipd'last_event, tpd_I1_O, TRUE),
                 2 => (I2_ipd'last_event, tpd_I2_O, TRUE),
                 3 => (I3_ipd'last_event, tpd_I3_O, TRUE),
                 4 => (I4_ipd'last_event, tpd_I4_O, TRUE),
                 5 => (I5_ipd'last_event, tpd_I5_O, TRUE),
                 6 => (I6_ipd'last_event, tpd_I6_O, TRUE),
                 7 => (I7_ipd'last_event, tpd_I7_O, TRUE),
                 8 => (I8_ipd'last_event, tpd_I8_O, TRUE),
                 9 => (I9_ipd'last_event, tpd_I9_O, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
 
end VITAL_VF;
 
configuration CFG_AND10_VITAL of AND10 is 
        for VITAL_VF
        end for; 
end CFG_AND10_VITAL;
----- VITAL model for cell AND11 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AND11 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_I0_O                       :	VitalDelayType01 := (3.050 ns, 3.050 ns);
      tpd_I1_O                       :	VitalDelayType01 := (3.050 ns, 3.050 ns);
      tpd_I2_O                       :	VitalDelayType01 := (3.050 ns, 3.050 ns);
      tpd_I3_O                       :	VitalDelayType01 := (3.050 ns, 3.050 ns);
      tpd_I4_O                       :	VitalDelayType01 := (3.050 ns, 3.050 ns);
      tpd_I5_O                       :	VitalDelayType01 := (3.050 ns, 3.050 ns);
      tpd_I6_O                       :	VitalDelayType01 := (3.050 ns, 3.050 ns);
      tpd_I7_O                       :	VitalDelayType01 := (3.050 ns, 3.050 ns);
      tpd_I8_O                       :	VitalDelayType01 := (3.050 ns, 3.050 ns);
      tpd_I9_O                       :	VitalDelayType01 := (3.050 ns, 3.050 ns);
      tpd_I10_O                      :	VitalDelayType01 := (3.050 ns, 3.050 ns);
      tipd_I0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I2                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I3                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I4                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I5                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I6                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I7                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I8                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I9                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I10                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      I0                             :	in    STD_ULOGIC;
      I1                             :	in    STD_ULOGIC;
      I2                             :	in    STD_ULOGIC;
      I3                             :	in    STD_ULOGIC;
      I4                             :	in    STD_ULOGIC;
      I5                             :	in    STD_ULOGIC;
      I6                             :	in    STD_ULOGIC;
      I7                             :	in    STD_ULOGIC;
      I8                             :	in    STD_ULOGIC;
      I9                             :	in    STD_ULOGIC;
      I10                            :	in    STD_ULOGIC;
      O                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AND11 : entity is TRUE;
end AND11;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
 
library VF1;
architecture VITAL_VF of AND11 is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL I0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I1_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I2_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I3_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I4_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I5_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I6_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I7_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I8_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I9_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I10_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (I0_ipd, I0, tipd_I0);
   VitalWireDelay (I1_ipd, I1, tipd_I1);
   VitalWireDelay (I2_ipd, I2, tipd_I2);
   VitalWireDelay (I3_ipd, I3, tipd_I3);
   VitalWireDelay (I4_ipd, I4, tipd_I4);
   VitalWireDelay (I5_ipd, I5, tipd_I5);
   VitalWireDelay (I6_ipd, I6, tipd_I6);
   VitalWireDelay (I7_ipd, I7, tipd_I7);
   VitalWireDelay (I8_ipd, I8, tipd_I8);
   VitalWireDelay (I9_ipd, I9, tipd_I9);
   VitalWireDelay (I10_ipd, I10, tipd_I10);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (I0_ipd, I1_ipd, I2_ipd, I3_ipd, I4_ipd, I5_ipd, I6_ipd, I7_ipd, I8_ipd, I9_ipd, I10_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS O_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE O_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      O_zd :=
       (I1_ipd) AND (I0_ipd) AND (I2_ipd) AND (I3_ipd) AND (I4_ipd) AND
         (I5_ipd) AND (I6_ipd) AND (I7_ipd) AND (I8_ipd) AND (I9_ipd) AND
         (I10_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => O,
       GlitchData => O_GlitchData,
       OutSignalName => "O",
       OutTemp => O_zd,
       Paths => (0 => (I0_ipd'last_event, tpd_I0_O, TRUE),
                 1 => (I1_ipd'last_event, tpd_I1_O, TRUE),
                 2 => (I2_ipd'last_event, tpd_I2_O, TRUE),
                 3 => (I3_ipd'last_event, tpd_I3_O, TRUE),
                 4 => (I4_ipd'last_event, tpd_I4_O, TRUE),
                 5 => (I5_ipd'last_event, tpd_I5_O, TRUE),
                 6 => (I6_ipd'last_event, tpd_I6_O, TRUE),
                 7 => (I7_ipd'last_event, tpd_I7_O, TRUE),
                 8 => (I8_ipd'last_event, tpd_I8_O, TRUE),
                 9 => (I9_ipd'last_event, tpd_I9_O, TRUE),
                 10 => (I10_ipd'last_event, tpd_I10_O, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;
 
configuration CFG_AND11_VITAL of AND11 is 
        for VITAL_VF
        end for; 
end CFG_AND11_VITAL;
----- VITAL model for cell AND12 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AND12 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_I0_O                       :	VitalDelayType01 := (3.050 ns, 3.050 ns);
      tpd_I1_O                       :	VitalDelayType01 := (3.050 ns, 3.050 ns);
      tpd_I2_O                       :	VitalDelayType01 := (3.050 ns, 3.050 ns);
      tpd_I3_O                       :	VitalDelayType01 := (3.050 ns, 3.050 ns);
      tpd_I4_O                       :	VitalDelayType01 := (3.050 ns, 3.050 ns);
      tpd_I5_O                       :	VitalDelayType01 := (3.050 ns, 3.050 ns);
      tpd_I6_O                       :	VitalDelayType01 := (3.050 ns, 3.050 ns);
      tpd_I7_O                       :	VitalDelayType01 := (3.050 ns, 3.050 ns);
      tpd_I8_O                       :	VitalDelayType01 := (3.050 ns, 3.050 ns);
      tpd_I9_O                       :	VitalDelayType01 := (3.050 ns, 3.050 ns);
      tpd_I10_O                      :	VitalDelayType01 := (3.050 ns, 3.050 ns);
      tpd_I11_O                      :	VitalDelayType01 := (3.050 ns, 3.050 ns);
      tipd_I0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I2                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I3                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I4                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I5                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I6                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I7                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I8                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I9                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I10                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I11                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      I0                             :	in    STD_ULOGIC;
      I1                             :	in    STD_ULOGIC;
      I2                             :	in    STD_ULOGIC;
      I3                             :	in    STD_ULOGIC;
      I4                             :	in    STD_ULOGIC;
      I5                             :	in    STD_ULOGIC;
      I6                             :	in    STD_ULOGIC;
      I7                             :	in    STD_ULOGIC;
      I8                             :	in    STD_ULOGIC;
      I9                             :	in    STD_ULOGIC;
      I10                            :	in    STD_ULOGIC;
      I11                            :	in    STD_ULOGIC;
      O                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AND12 : entity is TRUE;
end AND12;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
 
library VF1;
architecture VITAL_VF of AND12 is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL I0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I1_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I2_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I3_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I4_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I5_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I6_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I7_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I8_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I9_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I10_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I11_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (I0_ipd, I0, tipd_I0);
   VitalWireDelay (I1_ipd, I1, tipd_I1);
   VitalWireDelay (I2_ipd, I2, tipd_I2);
   VitalWireDelay (I3_ipd, I3, tipd_I3);
   VitalWireDelay (I4_ipd, I4, tipd_I4);
   VitalWireDelay (I5_ipd, I5, tipd_I5);
   VitalWireDelay (I6_ipd, I6, tipd_I6);
   VitalWireDelay (I7_ipd, I7, tipd_I7);
   VitalWireDelay (I8_ipd, I8, tipd_I8);
   VitalWireDelay (I9_ipd, I9, tipd_I9);
   VitalWireDelay (I10_ipd, I10, tipd_I10);
   VitalWireDelay (I11_ipd, I11, tipd_I11);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (I0_ipd, I1_ipd, I2_ipd, I3_ipd, I4_ipd, I5_ipd, I6_ipd, I7_ipd, I8_ipd, I9_ipd, I10_ipd, I11_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS O_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE O_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      O_zd :=
       (I1_ipd) AND (I0_ipd) AND (I2_ipd) AND (I3_ipd) AND (I4_ipd) AND
         (I5_ipd) AND (I6_ipd) AND (I7_ipd) AND (I8_ipd) AND (I9_ipd) AND
         (I10_ipd) AND (I11_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => O,
       GlitchData => O_GlitchData,
       OutSignalName => "O",
       OutTemp => O_zd,
       Paths => (0 => (I0_ipd'last_event, tpd_I0_O, TRUE),
                 1 => (I1_ipd'last_event, tpd_I1_O, TRUE),
                 2 => (I2_ipd'last_event, tpd_I2_O, TRUE),
                 3 => (I3_ipd'last_event, tpd_I3_O, TRUE),
                 4 => (I4_ipd'last_event, tpd_I4_O, TRUE),
                 5 => (I5_ipd'last_event, tpd_I5_O, TRUE),
                 6 => (I6_ipd'last_event, tpd_I6_O, TRUE),
                 7 => (I7_ipd'last_event, tpd_I7_O, TRUE),
                 8 => (I8_ipd'last_event, tpd_I8_O, TRUE),
                 9 => (I9_ipd'last_event, tpd_I9_O, TRUE),
                 10 => (I10_ipd'last_event, tpd_I10_O, TRUE),
                 11 => (I11_ipd'last_event, tpd_I11_O, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;
 
configuration CFG_AND12_VITAL of AND12 is 
        for VITAL_VF
        end for; 
end CFG_AND12_VITAL;
----- VITAL model for cell AND13 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AND13 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_I0_O                       :	VitalDelayType01 := (3.600 ns, 3.600 ns);
      tpd_I1_O                       :	VitalDelayType01 := (3.600 ns, 3.600 ns);
      tpd_I2_O                       :	VitalDelayType01 := (3.600 ns, 3.600 ns);
      tpd_I3_O                       :	VitalDelayType01 := (3.600 ns, 3.600 ns);
      tpd_I4_O                       :	VitalDelayType01 := (3.600 ns, 3.600 ns);
      tpd_I5_O                       :	VitalDelayType01 := (3.600 ns, 3.600 ns);
      tpd_I6_O                       :	VitalDelayType01 := (3.600 ns, 3.600 ns);
      tpd_I7_O                       :	VitalDelayType01 := (3.600 ns, 3.600 ns);
      tpd_I8_O                       :	VitalDelayType01 := (3.600 ns, 3.600 ns);
      tpd_I9_O                       :	VitalDelayType01 := (3.600 ns, 3.600 ns);
      tpd_I10_O                      :	VitalDelayType01 := (3.600 ns, 3.600 ns);
      tpd_I11_O                      :	VitalDelayType01 := (3.600 ns, 3.600 ns);
      tpd_I12_O                      :	VitalDelayType01 := (3.600 ns, 3.600 ns);
      tipd_I0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I2                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I3                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I4                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I5                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I6                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I7                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I8                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I9                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I10                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I11                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I12                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      I0                             :	in    STD_ULOGIC;
      I1                             :	in    STD_ULOGIC;
      I2                             :	in    STD_ULOGIC;
      I3                             :	in    STD_ULOGIC;
      I4                             :	in    STD_ULOGIC;
      I5                             :	in    STD_ULOGIC;
      I6                             :	in    STD_ULOGIC;
      I7                             :	in    STD_ULOGIC;
      I8                             :	in    STD_ULOGIC;
      I9                             :	in    STD_ULOGIC;
      I10                            :	in    STD_ULOGIC;
      I11                            :	in    STD_ULOGIC;
      I12                            :	in    STD_ULOGIC;
      O                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AND13 : entity is TRUE;
end AND13;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
 
library VF1;
architecture VITAL_VF of AND13 is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL I0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I1_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I2_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I3_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I4_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I5_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I6_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I7_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I8_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I9_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I10_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I11_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I12_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (I0_ipd, I0, tipd_I0);
   VitalWireDelay (I1_ipd, I1, tipd_I1);
   VitalWireDelay (I2_ipd, I2, tipd_I2);
   VitalWireDelay (I3_ipd, I3, tipd_I3);
   VitalWireDelay (I4_ipd, I4, tipd_I4);
   VitalWireDelay (I5_ipd, I5, tipd_I5);
   VitalWireDelay (I6_ipd, I6, tipd_I6);
   VitalWireDelay (I7_ipd, I7, tipd_I7);
   VitalWireDelay (I8_ipd, I8, tipd_I8);
   VitalWireDelay (I9_ipd, I9, tipd_I9);
   VitalWireDelay (I10_ipd, I10, tipd_I10);
   VitalWireDelay (I11_ipd, I11, tipd_I11);
   VitalWireDelay (I12_ipd, I12, tipd_I12);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (I0_ipd, I1_ipd, I2_ipd, I3_ipd, I4_ipd, I5_ipd, I6_ipd, I7_ipd, I8_ipd, I9_ipd, I10_ipd, I11_ipd, I12_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS O_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE O_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      O_zd :=
       (I1_ipd) AND (I0_ipd) AND (I2_ipd) AND (I3_ipd) AND (I4_ipd) AND
         (I5_ipd) AND (I6_ipd) AND (I7_ipd) AND (I8_ipd) AND (I9_ipd) AND
         (I10_ipd) AND (I11_ipd) AND (I12_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => O,
       GlitchData => O_GlitchData,
       OutSignalName => "O",
       OutTemp => O_zd,
       Paths => (0 => (I0_ipd'last_event, tpd_I0_O, TRUE),
                 1 => (I1_ipd'last_event, tpd_I1_O, TRUE),
                 2 => (I2_ipd'last_event, tpd_I2_O, TRUE),
                 3 => (I3_ipd'last_event, tpd_I3_O, TRUE),
                 4 => (I4_ipd'last_event, tpd_I4_O, TRUE),
                 5 => (I5_ipd'last_event, tpd_I5_O, TRUE),
                 6 => (I6_ipd'last_event, tpd_I6_O, TRUE),
                 7 => (I7_ipd'last_event, tpd_I7_O, TRUE),
                 8 => (I8_ipd'last_event, tpd_I8_O, TRUE),
                 9 => (I9_ipd'last_event, tpd_I9_O, TRUE),
                 10 => (I10_ipd'last_event, tpd_I10_O, TRUE),
                 11 => (I11_ipd'last_event, tpd_I11_O, TRUE),
                 12 => (I12_ipd'last_event, tpd_I12_O, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;
 
configuration CFG_AND13_VITAL of AND13 is 
        for VITAL_VF
        end for; 
end CFG_AND13_VITAL;
----- VITAL model for cell AND14 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AND14 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_I0_O                       :	VitalDelayType01 := (3.600 ns, 3.600 ns);
      tpd_I1_O                       :	VitalDelayType01 := (3.600 ns, 3.600 ns);
      tpd_I2_O                       :	VitalDelayType01 := (3.600 ns, 3.600 ns);
      tpd_I3_O                       :	VitalDelayType01 := (3.600 ns, 3.600 ns);
      tpd_I4_O                       :	VitalDelayType01 := (3.600 ns, 3.600 ns);
      tpd_I5_O                       :	VitalDelayType01 := (3.600 ns, 3.600 ns);
      tpd_I6_O                       :	VitalDelayType01 := (3.600 ns, 3.600 ns);
      tpd_I7_O                       :	VitalDelayType01 := (3.600 ns, 3.600 ns);
      tpd_I8_O                       :	VitalDelayType01 := (3.600 ns, 3.600 ns);
      tpd_I9_O                       :	VitalDelayType01 := (3.600 ns, 3.600 ns);
      tpd_I10_O                      :	VitalDelayType01 := (3.600 ns, 3.600 ns);
      tpd_I11_O                      :	VitalDelayType01 := (3.600 ns, 3.600 ns);
      tpd_I12_O                      :	VitalDelayType01 := (3.600 ns, 3.600 ns);
      tpd_I13_O                      :	VitalDelayType01 := (3.600 ns, 3.600 ns);
      tipd_I0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I2                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I3                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I4                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I5                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I6                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I7                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I8                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I9                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I10                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I11                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I12                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I13                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      I0                             :	in    STD_ULOGIC;
      I1                             :	in    STD_ULOGIC;
      I2                             :	in    STD_ULOGIC;
      I3                             :	in    STD_ULOGIC;
      I4                             :	in    STD_ULOGIC;
      I5                             :	in    STD_ULOGIC;
      I6                             :	in    STD_ULOGIC;
      I7                             :	in    STD_ULOGIC;
      I8                             :	in    STD_ULOGIC;
      I9                             :	in    STD_ULOGIC;
      I10                            :	in    STD_ULOGIC;
      I11                            :	in    STD_ULOGIC;
      I12                            :	in    STD_ULOGIC;
      I13                            :	in    STD_ULOGIC;
      O                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AND14 : entity is TRUE;
end AND14;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
 
library VF1;
architecture VITAL_VF of AND14 is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL I0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I1_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I2_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I3_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I4_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I5_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I6_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I7_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I8_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I9_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I10_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I11_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I12_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I13_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (I0_ipd, I0, tipd_I0);
   VitalWireDelay (I1_ipd, I1, tipd_I1);
   VitalWireDelay (I2_ipd, I2, tipd_I2);
   VitalWireDelay (I3_ipd, I3, tipd_I3);
   VitalWireDelay (I4_ipd, I4, tipd_I4);
   VitalWireDelay (I5_ipd, I5, tipd_I5);
   VitalWireDelay (I6_ipd, I6, tipd_I6);
   VitalWireDelay (I7_ipd, I7, tipd_I7);
   VitalWireDelay (I8_ipd, I8, tipd_I8);
   VitalWireDelay (I9_ipd, I9, tipd_I9);
   VitalWireDelay (I10_ipd, I10, tipd_I10);
   VitalWireDelay (I11_ipd, I11, tipd_I11);
   VitalWireDelay (I12_ipd, I12, tipd_I12);
   VitalWireDelay (I13_ipd, I13, tipd_I13);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (I0_ipd, I1_ipd, I2_ipd, I3_ipd, I4_ipd, I5_ipd, I6_ipd, I7_ipd, I8_ipd, I9_ipd, I10_ipd, I11_ipd, I12_ipd, I13_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS O_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE O_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      O_zd :=
       (I1_ipd) AND (I0_ipd) AND (I2_ipd) AND (I3_ipd) AND (I4_ipd) AND
         (I5_ipd) AND (I6_ipd) AND (I7_ipd) AND (I8_ipd) AND (I9_ipd) AND
         (I10_ipd) AND (I11_ipd) AND (I12_ipd) AND (I13_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => O,
       GlitchData => O_GlitchData,
       OutSignalName => "O",
       OutTemp => O_zd,
       Paths => (0 => (I0_ipd'last_event, tpd_I0_O, TRUE),
                 1 => (I1_ipd'last_event, tpd_I1_O, TRUE),
                 2 => (I2_ipd'last_event, tpd_I2_O, TRUE),
                 3 => (I3_ipd'last_event, tpd_I3_O, TRUE),
                 4 => (I4_ipd'last_event, tpd_I4_O, TRUE),
                 5 => (I5_ipd'last_event, tpd_I5_O, TRUE),
                 6 => (I6_ipd'last_event, tpd_I6_O, TRUE),
                 7 => (I7_ipd'last_event, tpd_I7_O, TRUE),
                 8 => (I8_ipd'last_event, tpd_I8_O, TRUE),
                 9 => (I9_ipd'last_event, tpd_I9_O, TRUE),
                 10 => (I10_ipd'last_event, tpd_I10_O, TRUE),
                 11 => (I11_ipd'last_event, tpd_I11_O, TRUE),
                 12 => (I12_ipd'last_event, tpd_I12_O, TRUE),
                 13 => (I13_ipd'last_event, tpd_I13_O, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;
 
configuration CFG_AND14_VITAL of AND14 is 
        for VITAL_VF
        end for; 
end CFG_AND14_VITAL;
----- VITAL model for cell AND15 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AND15 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_I0_O                       :	VitalDelayType01 := (3.600 ns, 3.600 ns);
      tpd_I1_O                       :	VitalDelayType01 := (3.600 ns, 3.600 ns);
      tpd_I2_O                       :	VitalDelayType01 := (3.600 ns, 3.600 ns);
      tpd_I3_O                       :	VitalDelayType01 := (3.600 ns, 3.600 ns);
      tpd_I4_O                       :	VitalDelayType01 := (3.600 ns, 3.600 ns);
      tpd_I5_O                       :	VitalDelayType01 := (3.600 ns, 3.600 ns);
      tpd_I6_O                       :	VitalDelayType01 := (3.600 ns, 3.600 ns);
      tpd_I7_O                       :	VitalDelayType01 := (3.600 ns, 3.600 ns);
      tpd_I8_O                       :	VitalDelayType01 := (3.600 ns, 3.600 ns);
      tpd_I9_O                       :	VitalDelayType01 := (3.600 ns, 3.600 ns);
      tpd_I10_O                      :	VitalDelayType01 := (3.600 ns, 3.600 ns);
      tpd_I11_O                      :	VitalDelayType01 := (3.600 ns, 3.600 ns);
      tpd_I12_O                      :	VitalDelayType01 := (3.600 ns, 3.600 ns);
      tpd_I13_O                      :	VitalDelayType01 := (3.600 ns, 3.600 ns);
      tpd_I14_O                      :	VitalDelayType01 := (3.600 ns, 3.600 ns);
      tipd_I0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I2                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I3                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I4                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I5                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I6                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I7                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I8                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I9                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I10                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I11                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I12                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I13                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I14                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      I0                             :	in    STD_ULOGIC;
      I1                             :	in    STD_ULOGIC;
      I2                             :	in    STD_ULOGIC;
      I3                             :	in    STD_ULOGIC;
      I4                             :	in    STD_ULOGIC;
      I5                             :	in    STD_ULOGIC;
      I6                             :	in    STD_ULOGIC;
      I7                             :	in    STD_ULOGIC;
      I8                             :	in    STD_ULOGIC;
      I9                             :	in    STD_ULOGIC;
      I10                            :	in    STD_ULOGIC;
      I11                            :	in    STD_ULOGIC;
      I12                            :	in    STD_ULOGIC;
      I13                            :	in    STD_ULOGIC;
      I14                            :	in    STD_ULOGIC;
      O                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AND15 : entity is TRUE;
end AND15;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
 
library VF1;
architecture VITAL_VF of AND15 is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL I0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I1_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I2_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I3_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I4_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I5_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I6_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I7_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I8_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I9_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I10_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I11_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I12_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I13_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I14_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (I0_ipd, I0, tipd_I0);
   VitalWireDelay (I1_ipd, I1, tipd_I1);
   VitalWireDelay (I2_ipd, I2, tipd_I2);
   VitalWireDelay (I3_ipd, I3, tipd_I3);
   VitalWireDelay (I4_ipd, I4, tipd_I4);
   VitalWireDelay (I5_ipd, I5, tipd_I5);
   VitalWireDelay (I6_ipd, I6, tipd_I6);
   VitalWireDelay (I7_ipd, I7, tipd_I7);
   VitalWireDelay (I8_ipd, I8, tipd_I8);
   VitalWireDelay (I9_ipd, I9, tipd_I9);
   VitalWireDelay (I10_ipd, I10, tipd_I10);
   VitalWireDelay (I11_ipd, I11, tipd_I11);
   VitalWireDelay (I12_ipd, I12, tipd_I12);
   VitalWireDelay (I13_ipd, I13, tipd_I13);
   VitalWireDelay (I14_ipd, I14, tipd_I14);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (I0_ipd, I1_ipd, I2_ipd, I3_ipd, I4_ipd, I5_ipd, I6_ipd, I7_ipd, I8_ipd, I9_ipd, I10_ipd, I11_ipd, I12_ipd, I13_ipd, I14_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS O_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE O_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      O_zd :=
       (I1_ipd) AND (I0_ipd) AND (I2_ipd) AND (I3_ipd) AND (I4_ipd) AND
         (I5_ipd) AND (I6_ipd) AND (I7_ipd) AND (I8_ipd) AND (I9_ipd) AND
         (I10_ipd) AND (I11_ipd) AND (I12_ipd) AND (I13_ipd) AND (I14_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => O,
       GlitchData => O_GlitchData,
       OutSignalName => "O",
       OutTemp => O_zd,
       Paths => (0 => (I0_ipd'last_event, tpd_I0_O, TRUE),
                 1 => (I1_ipd'last_event, tpd_I1_O, TRUE),
                 2 => (I2_ipd'last_event, tpd_I2_O, TRUE),
                 3 => (I3_ipd'last_event, tpd_I3_O, TRUE),
                 4 => (I4_ipd'last_event, tpd_I4_O, TRUE),
                 5 => (I5_ipd'last_event, tpd_I5_O, TRUE),
                 6 => (I6_ipd'last_event, tpd_I6_O, TRUE),
                 7 => (I7_ipd'last_event, tpd_I7_O, TRUE),
                 8 => (I8_ipd'last_event, tpd_I8_O, TRUE),
                 9 => (I9_ipd'last_event, tpd_I9_O, TRUE),
                 10 => (I10_ipd'last_event, tpd_I10_O, TRUE),
                 11 => (I11_ipd'last_event, tpd_I11_O, TRUE),
                 12 => (I12_ipd'last_event, tpd_I12_O, TRUE),
                 13 => (I13_ipd'last_event, tpd_I13_O, TRUE),
                 14 => (I14_ipd'last_event, tpd_I14_O, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;
 
configuration CFG_AND15_VITAL of AND15 is 
        for VITAL_VF
        end for; 
end CFG_AND15_VITAL;
----- VITAL model for cell AND16 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AND16 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_I0_O                       :	VitalDelayType01 := (3.600 ns, 3.600 ns);
      tpd_I1_O                       :	VitalDelayType01 := (3.600 ns, 3.600 ns);
      tpd_I2_O                       :	VitalDelayType01 := (3.600 ns, 3.600 ns);
      tpd_I3_O                       :	VitalDelayType01 := (3.600 ns, 3.600 ns);
      tpd_I4_O                       :	VitalDelayType01 := (3.600 ns, 3.600 ns);
      tpd_I5_O                       :	VitalDelayType01 := (3.600 ns, 3.600 ns);
      tpd_I6_O                       :	VitalDelayType01 := (3.600 ns, 3.600 ns);
      tpd_I7_O                       :	VitalDelayType01 := (3.600 ns, 3.600 ns);
      tpd_I8_O                       :	VitalDelayType01 := (3.600 ns, 3.600 ns);
      tpd_I9_O                       :	VitalDelayType01 := (3.600 ns, 3.600 ns);
      tpd_I10_O                      :	VitalDelayType01 := (3.600 ns, 3.600 ns);
      tpd_I11_O                      :	VitalDelayType01 := (3.600 ns, 3.600 ns);
      tpd_I12_O                      :	VitalDelayType01 := (3.600 ns, 3.600 ns);
      tpd_I13_O                      :	VitalDelayType01 := (3.600 ns, 3.600 ns);
      tpd_I14_O                      :	VitalDelayType01 := (3.600 ns, 3.600 ns);
      tpd_I15_O                      :	VitalDelayType01 := (3.600 ns, 3.600 ns);
      tipd_I0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I2                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I3                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I4                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I5                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I6                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I7                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I8                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I9                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I10                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I11                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I12                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I13                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I14                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I15                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      I0                             :	in    STD_ULOGIC;
      I1                             :	in    STD_ULOGIC;
      I2                             :	in    STD_ULOGIC;
      I3                             :	in    STD_ULOGIC;
      I4                             :	in    STD_ULOGIC;
      I5                             :	in    STD_ULOGIC;
      I6                             :	in    STD_ULOGIC;
      I7                             :	in    STD_ULOGIC;
      I8                             :	in    STD_ULOGIC;
      I9                             :	in    STD_ULOGIC;
      I10                            :	in    STD_ULOGIC;
      I11                            :	in    STD_ULOGIC;
      I12                            :	in    STD_ULOGIC;
      I13                            :	in    STD_ULOGIC;
      I14                            :	in    STD_ULOGIC;
      I15                            :	in    STD_ULOGIC;
      O                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AND16 : entity is TRUE;
end AND16;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
 
library VF1;
architecture VITAL_VF of AND16 is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL I0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I1_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I2_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I3_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I4_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I5_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I6_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I7_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I8_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I9_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I10_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I11_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I12_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I13_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I14_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I15_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (I0_ipd, I0, tipd_I0);
   VitalWireDelay (I1_ipd, I1, tipd_I1);
   VitalWireDelay (I2_ipd, I2, tipd_I2);
   VitalWireDelay (I3_ipd, I3, tipd_I3);
   VitalWireDelay (I4_ipd, I4, tipd_I4);
   VitalWireDelay (I5_ipd, I5, tipd_I5);
   VitalWireDelay (I6_ipd, I6, tipd_I6);
   VitalWireDelay (I7_ipd, I7, tipd_I7);
   VitalWireDelay (I8_ipd, I8, tipd_I8);
   VitalWireDelay (I9_ipd, I9, tipd_I9);
   VitalWireDelay (I10_ipd, I10, tipd_I10);
   VitalWireDelay (I11_ipd, I11, tipd_I11);
   VitalWireDelay (I12_ipd, I12, tipd_I12);
   VitalWireDelay (I13_ipd, I13, tipd_I13);
   VitalWireDelay (I14_ipd, I14, tipd_I14);
   VitalWireDelay (I15_ipd, I15, tipd_I15);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (I0_ipd, I1_ipd, I2_ipd, I3_ipd, I4_ipd, I5_ipd, I6_ipd, I7_ipd, I8_ipd, I9_ipd, I10_ipd, I11_ipd, I12_ipd, I13_ipd, I14_ipd, I15_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS O_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE O_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      O_zd :=
       (I1_ipd) AND (I0_ipd) AND (I2_ipd) AND (I3_ipd) AND (I4_ipd) AND
         (I5_ipd) AND (I6_ipd) AND (I7_ipd) AND (I8_ipd) AND (I9_ipd) AND
         (I10_ipd) AND (I11_ipd) AND (I12_ipd) AND (I13_ipd) AND (I14_ipd)
         AND (I15_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => O,
       GlitchData => O_GlitchData,
       OutSignalName => "O",
       OutTemp => O_zd,
       Paths => (0 => (I0_ipd'last_event, tpd_I0_O, TRUE),
                 1 => (I1_ipd'last_event, tpd_I1_O, TRUE),
                 2 => (I2_ipd'last_event, tpd_I2_O, TRUE),
                 3 => (I3_ipd'last_event, tpd_I3_O, TRUE),
                 4 => (I4_ipd'last_event, tpd_I4_O, TRUE),
                 5 => (I5_ipd'last_event, tpd_I5_O, TRUE),
                 6 => (I6_ipd'last_event, tpd_I6_O, TRUE),
                 7 => (I7_ipd'last_event, tpd_I7_O, TRUE),
                 8 => (I8_ipd'last_event, tpd_I8_O, TRUE),
                 9 => (I9_ipd'last_event, tpd_I9_O, TRUE),
                 10 => (I10_ipd'last_event, tpd_I10_O, TRUE),
                 11 => (I11_ipd'last_event, tpd_I11_O, TRUE),
                 12 => (I12_ipd'last_event, tpd_I12_O, TRUE),
                 13 => (I13_ipd'last_event, tpd_I13_O, TRUE),
                 14 => (I14_ipd'last_event, tpd_I14_O, TRUE),
                 15 => (I15_ipd'last_event, tpd_I15_O, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;
 
configuration CFG_AND16_VITAL of AND16 is 
        for VITAL_VF
        end for; 
end CFG_AND16_VITAL;
----- VITAL model for cell AND17 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AND17 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_I0_O                       :	VitalDelayType01 := (4.300 ns, 4.300 ns);
      tpd_I1_O                       :	VitalDelayType01 := (4.300 ns, 4.300 ns);
      tpd_I2_O                       :	VitalDelayType01 := (4.300 ns, 4.300 ns);
      tpd_I3_O                       :	VitalDelayType01 := (4.300 ns, 4.300 ns);
      tpd_I4_O                       :	VitalDelayType01 := (4.300 ns, 4.300 ns);
      tpd_I5_O                       :	VitalDelayType01 := (4.300 ns, 4.300 ns);
      tpd_I6_O                       :	VitalDelayType01 := (4.300 ns, 4.300 ns);
      tpd_I7_O                       :	VitalDelayType01 := (4.300 ns, 4.300 ns);
      tpd_I8_O                       :	VitalDelayType01 := (4.300 ns, 4.300 ns);
      tpd_I9_O                       :	VitalDelayType01 := (4.300 ns, 4.300 ns);
      tpd_I10_O                      :	VitalDelayType01 := (4.300 ns, 4.300 ns);
      tpd_I11_O                      :	VitalDelayType01 := (4.300 ns, 4.300 ns);
      tpd_I12_O                      :	VitalDelayType01 := (4.300 ns, 4.300 ns);
      tpd_I13_O                      :	VitalDelayType01 := (4.300 ns, 4.300 ns);
      tpd_I14_O                      :	VitalDelayType01 := (4.300 ns, 4.300 ns);
      tpd_I15_O                      :	VitalDelayType01 := (4.300 ns, 4.300 ns);
      tpd_I16_O                      :	VitalDelayType01 := (4.300 ns, 4.300 ns);
      tipd_I0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I2                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I3                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I4                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I5                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I6                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I7                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I8                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I9                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I10                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I11                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I12                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I13                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I14                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I15                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I16                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      I0                             :	in    STD_ULOGIC;
      I1                             :	in    STD_ULOGIC;
      I2                             :	in    STD_ULOGIC;
      I3                             :	in    STD_ULOGIC;
      I4                             :	in    STD_ULOGIC;
      I5                             :	in    STD_ULOGIC;
      I6                             :	in    STD_ULOGIC;
      I7                             :	in    STD_ULOGIC;
      I8                             :	in    STD_ULOGIC;
      I9                             :	in    STD_ULOGIC;
      I10                            :	in    STD_ULOGIC;
      I11                            :	in    STD_ULOGIC;
      I12                            :	in    STD_ULOGIC;
      I13                            :	in    STD_ULOGIC;
      I14                            :	in    STD_ULOGIC;
      I15                            :	in    STD_ULOGIC;
      I16                            :	in    STD_ULOGIC;
      O                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AND17 : entity is TRUE;
end AND17;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
 
library VF1;
architecture VITAL_VF of AND17 is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL I0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I1_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I2_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I3_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I4_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I5_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I6_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I7_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I8_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I9_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I10_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I11_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I12_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I13_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I14_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I15_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I16_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (I0_ipd, I0, tipd_I0);
   VitalWireDelay (I1_ipd, I1, tipd_I1);
   VitalWireDelay (I2_ipd, I2, tipd_I2);
   VitalWireDelay (I3_ipd, I3, tipd_I3);
   VitalWireDelay (I4_ipd, I4, tipd_I4);
   VitalWireDelay (I5_ipd, I5, tipd_I5);
   VitalWireDelay (I6_ipd, I6, tipd_I6);
   VitalWireDelay (I7_ipd, I7, tipd_I7);
   VitalWireDelay (I8_ipd, I8, tipd_I8);
   VitalWireDelay (I9_ipd, I9, tipd_I9);
   VitalWireDelay (I10_ipd, I10, tipd_I10);
   VitalWireDelay (I11_ipd, I11, tipd_I11);
   VitalWireDelay (I12_ipd, I12, tipd_I12);
   VitalWireDelay (I13_ipd, I13, tipd_I13);
   VitalWireDelay (I14_ipd, I14, tipd_I14);
   VitalWireDelay (I15_ipd, I15, tipd_I15);
   VitalWireDelay (I16_ipd, I16, tipd_I16);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (I0_ipd, I1_ipd, I2_ipd, I3_ipd, I4_ipd, I5_ipd, I6_ipd, I7_ipd, I8_ipd, I9_ipd, I10_ipd, I11_ipd, I12_ipd, I13_ipd, I14_ipd, I15_ipd, I16_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS O_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE O_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      O_zd :=
       (I1_ipd) AND (I0_ipd) AND (I2_ipd) AND (I3_ipd) AND (I4_ipd) AND
         (I5_ipd) AND (I6_ipd) AND (I7_ipd) AND (I8_ipd) AND (I9_ipd) AND
         (I10_ipd) AND (I11_ipd) AND (I12_ipd) AND (I13_ipd) AND (I14_ipd)
         AND (I15_ipd) AND (I16_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => O,
       GlitchData => O_GlitchData,
       OutSignalName => "O",
       OutTemp => O_zd,
       Paths => (0 => (I0_ipd'last_event, tpd_I0_O, TRUE),
                 1 => (I1_ipd'last_event, tpd_I1_O, TRUE),
                 2 => (I2_ipd'last_event, tpd_I2_O, TRUE),
                 3 => (I3_ipd'last_event, tpd_I3_O, TRUE),
                 4 => (I4_ipd'last_event, tpd_I4_O, TRUE),
                 5 => (I5_ipd'last_event, tpd_I5_O, TRUE),
                 6 => (I6_ipd'last_event, tpd_I6_O, TRUE),
                 7 => (I7_ipd'last_event, tpd_I7_O, TRUE),
                 8 => (I8_ipd'last_event, tpd_I8_O, TRUE),
                 9 => (I9_ipd'last_event, tpd_I9_O, TRUE),
                 10 => (I10_ipd'last_event, tpd_I10_O, TRUE),
                 11 => (I11_ipd'last_event, tpd_I11_O, TRUE),
                 12 => (I12_ipd'last_event, tpd_I12_O, TRUE),
                 13 => (I13_ipd'last_event, tpd_I13_O, TRUE),
                 14 => (I14_ipd'last_event, tpd_I14_O, TRUE),
                 15 => (I15_ipd'last_event, tpd_I15_O, TRUE),
                 16 => (I16_ipd'last_event, tpd_I16_O, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;
 
configuration CFG_AND17_VITAL of AND17 is 
        for VITAL_VF
        end for; 
end CFG_AND17_VITAL;
----- VITAL model for cell AND18 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AND18 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_I0_O                       :	VitalDelayType01 := (4.300 ns, 4.300 ns);
      tpd_I1_O                       :	VitalDelayType01 := (4.300 ns, 4.300 ns);
      tpd_I2_O                       :	VitalDelayType01 := (4.300 ns, 4.300 ns);
      tpd_I3_O                       :	VitalDelayType01 := (4.300 ns, 4.300 ns);
      tpd_I4_O                       :	VitalDelayType01 := (4.300 ns, 4.300 ns);
      tpd_I5_O                       :	VitalDelayType01 := (4.300 ns, 4.300 ns);
      tpd_I6_O                       :	VitalDelayType01 := (4.300 ns, 4.300 ns);
      tpd_I7_O                       :	VitalDelayType01 := (4.300 ns, 4.300 ns);
      tpd_I8_O                       :	VitalDelayType01 := (4.300 ns, 4.300 ns);
      tpd_I9_O                       :	VitalDelayType01 := (4.300 ns, 4.300 ns);
      tpd_I10_O                      :	VitalDelayType01 := (4.300 ns, 4.300 ns);
      tpd_I11_O                      :	VitalDelayType01 := (4.300 ns, 4.300 ns);
      tpd_I12_O                      :	VitalDelayType01 := (4.300 ns, 4.300 ns);
      tpd_I13_O                      :	VitalDelayType01 := (4.300 ns, 4.300 ns);
      tpd_I14_O                      :	VitalDelayType01 := (4.300 ns, 4.300 ns);
      tpd_I15_O                      :	VitalDelayType01 := (4.300 ns, 4.300 ns);
      tpd_I16_O                      :	VitalDelayType01 := (4.300 ns, 4.300 ns);
      tpd_I17_O                      :	VitalDelayType01 := (4.300 ns, 4.300 ns);
      tipd_I0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I2                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I3                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I4                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I5                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I6                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I7                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I8                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I9                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I10                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I11                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I12                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I13                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I14                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I15                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I16                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I17                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      I0                             :	in    STD_ULOGIC;
      I1                             :	in    STD_ULOGIC;
      I2                             :	in    STD_ULOGIC;
      I3                             :	in    STD_ULOGIC;
      I4                             :	in    STD_ULOGIC;
      I5                             :	in    STD_ULOGIC;
      I6                             :	in    STD_ULOGIC;
      I7                             :	in    STD_ULOGIC;
      I8                             :	in    STD_ULOGIC;
      I9                             :	in    STD_ULOGIC;
      I10                            :	in    STD_ULOGIC;
      I11                            :	in    STD_ULOGIC;
      I12                            :	in    STD_ULOGIC;
      I13                            :	in    STD_ULOGIC;
      I14                            :	in    STD_ULOGIC;
      I15                            :	in    STD_ULOGIC;
      I16                            :	in    STD_ULOGIC;
      I17                            :	in    STD_ULOGIC;
      O                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AND18 : entity is TRUE;
end AND18;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
 
library VF1;
architecture VITAL_VF of AND18 is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL I0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I1_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I2_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I3_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I4_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I5_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I6_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I7_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I8_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I9_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I10_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I11_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I12_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I13_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I14_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I15_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I16_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I17_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (I0_ipd, I0, tipd_I0);
   VitalWireDelay (I1_ipd, I1, tipd_I1);
   VitalWireDelay (I2_ipd, I2, tipd_I2);
   VitalWireDelay (I3_ipd, I3, tipd_I3);
   VitalWireDelay (I4_ipd, I4, tipd_I4);
   VitalWireDelay (I5_ipd, I5, tipd_I5);
   VitalWireDelay (I6_ipd, I6, tipd_I6);
   VitalWireDelay (I7_ipd, I7, tipd_I7);
   VitalWireDelay (I8_ipd, I8, tipd_I8);
   VitalWireDelay (I9_ipd, I9, tipd_I9);
   VitalWireDelay (I10_ipd, I10, tipd_I10);
   VitalWireDelay (I11_ipd, I11, tipd_I11);
   VitalWireDelay (I12_ipd, I12, tipd_I12);
   VitalWireDelay (I13_ipd, I13, tipd_I13);
   VitalWireDelay (I14_ipd, I14, tipd_I14);
   VitalWireDelay (I15_ipd, I15, tipd_I15);
   VitalWireDelay (I16_ipd, I16, tipd_I16);
   VitalWireDelay (I17_ipd, I17, tipd_I17);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (I0_ipd, I1_ipd, I2_ipd, I3_ipd, I4_ipd, I5_ipd, I6_ipd, I7_ipd, I8_ipd, I9_ipd, I10_ipd, I11_ipd, I12_ipd, I13_ipd, I14_ipd, I15_ipd, I16_ipd, I17_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS O_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE O_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      O_zd :=
       (I1_ipd) AND (I0_ipd) AND (I2_ipd) AND (I3_ipd) AND (I4_ipd) AND
         (I5_ipd) AND (I6_ipd) AND (I7_ipd) AND (I8_ipd) AND (I9_ipd) AND
         (I10_ipd) AND (I11_ipd) AND (I12_ipd) AND (I13_ipd) AND (I14_ipd)
         AND (I15_ipd) AND (I16_ipd) AND (I17_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => O,
       GlitchData => O_GlitchData,
       OutSignalName => "O",
       OutTemp => O_zd,
       Paths => (0 => (I0_ipd'last_event, tpd_I0_O, TRUE),
                 1 => (I1_ipd'last_event, tpd_I1_O, TRUE),
                 2 => (I2_ipd'last_event, tpd_I2_O, TRUE),
                 3 => (I3_ipd'last_event, tpd_I3_O, TRUE),
                 4 => (I4_ipd'last_event, tpd_I4_O, TRUE),
                 5 => (I5_ipd'last_event, tpd_I5_O, TRUE),
                 6 => (I6_ipd'last_event, tpd_I6_O, TRUE),
                 7 => (I7_ipd'last_event, tpd_I7_O, TRUE),
                 8 => (I8_ipd'last_event, tpd_I8_O, TRUE),
                 9 => (I9_ipd'last_event, tpd_I9_O, TRUE),
                 10 => (I10_ipd'last_event, tpd_I10_O, TRUE),
                 11 => (I11_ipd'last_event, tpd_I11_O, TRUE),
                 12 => (I12_ipd'last_event, tpd_I12_O, TRUE),
                 13 => (I13_ipd'last_event, tpd_I13_O, TRUE),
                 14 => (I14_ipd'last_event, tpd_I14_O, TRUE),
                 15 => (I15_ipd'last_event, tpd_I15_O, TRUE),
                 16 => (I16_ipd'last_event, tpd_I16_O, TRUE),
                 17 => (I17_ipd'last_event, tpd_I17_O, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;
 
configuration CFG_AND18_VITAL of AND18 is 
        for VITAL_VF
        end for; 
end CFG_AND18_VITAL;
----- VITAL model for cell AND19 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AND19 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_I0_O                       :	VitalDelayType01 := (4.300 ns, 4.300 ns);
      tpd_I1_O                       :	VitalDelayType01 := (4.300 ns, 4.300 ns);
      tpd_I2_O                       :	VitalDelayType01 := (4.300 ns, 4.300 ns);
      tpd_I3_O                       :	VitalDelayType01 := (4.300 ns, 4.300 ns);
      tpd_I4_O                       :	VitalDelayType01 := (4.300 ns, 4.300 ns);
      tpd_I5_O                       :	VitalDelayType01 := (4.300 ns, 4.300 ns);
      tpd_I6_O                       :	VitalDelayType01 := (4.300 ns, 4.300 ns);
      tpd_I7_O                       :	VitalDelayType01 := (4.300 ns, 4.300 ns);
      tpd_I8_O                       :	VitalDelayType01 := (4.300 ns, 4.300 ns);
      tpd_I9_O                       :	VitalDelayType01 := (4.300 ns, 4.300 ns);
      tpd_I10_O                      :	VitalDelayType01 := (4.300 ns, 4.300 ns);
      tpd_I11_O                      :	VitalDelayType01 := (4.300 ns, 4.300 ns);
      tpd_I12_O                      :	VitalDelayType01 := (4.300 ns, 4.300 ns);
      tpd_I13_O                      :	VitalDelayType01 := (4.300 ns, 4.300 ns);
      tpd_I14_O                      :	VitalDelayType01 := (4.300 ns, 4.300 ns);
      tpd_I15_O                      :	VitalDelayType01 := (4.300 ns, 4.300 ns);
      tpd_I16_O                      :	VitalDelayType01 := (4.300 ns, 4.300 ns);
      tpd_I17_O                      :	VitalDelayType01 := (4.300 ns, 4.300 ns);
      tpd_I18_O                      :	VitalDelayType01 := (4.300 ns, 4.300 ns);
      tipd_I0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I2                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I3                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I4                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I5                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I6                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I7                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I8                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I9                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I10                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I11                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I12                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I13                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I14                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I15                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I16                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I17                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I18                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      I0                             :	in    STD_ULOGIC;
      I1                             :	in    STD_ULOGIC;
      I2                             :	in    STD_ULOGIC;
      I3                             :	in    STD_ULOGIC;
      I4                             :	in    STD_ULOGIC;
      I5                             :	in    STD_ULOGIC;
      I6                             :	in    STD_ULOGIC;
      I7                             :	in    STD_ULOGIC;
      I8                             :	in    STD_ULOGIC;
      I9                             :	in    STD_ULOGIC;
      I10                            :	in    STD_ULOGIC;
      I11                            :	in    STD_ULOGIC;
      I12                            :	in    STD_ULOGIC;
      I13                            :	in    STD_ULOGIC;
      I14                            :	in    STD_ULOGIC;
      I15                            :	in    STD_ULOGIC;
      I16                            :	in    STD_ULOGIC;
      I17                            :	in    STD_ULOGIC;
      I18                            :	in    STD_ULOGIC;
      O                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AND19 : entity is TRUE;
end AND19;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
 
library VF1;
architecture VITAL_VF of AND19 is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL I0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I1_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I2_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I3_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I4_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I5_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I6_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I7_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I8_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I9_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I10_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I11_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I12_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I13_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I14_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I15_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I16_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I17_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I18_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (I0_ipd, I0, tipd_I0);
   VitalWireDelay (I1_ipd, I1, tipd_I1);
   VitalWireDelay (I2_ipd, I2, tipd_I2);
   VitalWireDelay (I3_ipd, I3, tipd_I3);
   VitalWireDelay (I4_ipd, I4, tipd_I4);
   VitalWireDelay (I5_ipd, I5, tipd_I5);
   VitalWireDelay (I6_ipd, I6, tipd_I6);
   VitalWireDelay (I7_ipd, I7, tipd_I7);
   VitalWireDelay (I8_ipd, I8, tipd_I8);
   VitalWireDelay (I9_ipd, I9, tipd_I9);
   VitalWireDelay (I10_ipd, I10, tipd_I10);
   VitalWireDelay (I11_ipd, I11, tipd_I11);
   VitalWireDelay (I12_ipd, I12, tipd_I12);
   VitalWireDelay (I13_ipd, I13, tipd_I13);
   VitalWireDelay (I14_ipd, I14, tipd_I14);
   VitalWireDelay (I15_ipd, I15, tipd_I15);
   VitalWireDelay (I16_ipd, I16, tipd_I16);
   VitalWireDelay (I17_ipd, I17, tipd_I17);
   VitalWireDelay (I18_ipd, I18, tipd_I18);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (I0_ipd, I1_ipd, I2_ipd, I3_ipd, I4_ipd, I5_ipd, I6_ipd, I7_ipd, I8_ipd, I9_ipd, I10_ipd, I11_ipd, I12_ipd, I13_ipd, I14_ipd, I15_ipd, I16_ipd, I17_ipd, I18_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS O_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE O_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      O_zd :=
       (I1_ipd) AND (I0_ipd) AND (I2_ipd) AND (I3_ipd) AND (I4_ipd) AND
         (I5_ipd) AND (I6_ipd) AND (I7_ipd) AND (I8_ipd) AND (I9_ipd) AND
         (I10_ipd) AND (I11_ipd) AND (I12_ipd) AND (I13_ipd) AND (I14_ipd)
         AND (I15_ipd) AND (I16_ipd) AND (I17_ipd) AND (I18_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => O,
       GlitchData => O_GlitchData,
       OutSignalName => "O",
       OutTemp => O_zd,
       Paths => (0 => (I0_ipd'last_event, tpd_I0_O, TRUE),
                 1 => (I1_ipd'last_event, tpd_I1_O, TRUE),
                 2 => (I2_ipd'last_event, tpd_I2_O, TRUE),
                 3 => (I3_ipd'last_event, tpd_I3_O, TRUE),
                 4 => (I4_ipd'last_event, tpd_I4_O, TRUE),
                 5 => (I5_ipd'last_event, tpd_I5_O, TRUE),
                 6 => (I6_ipd'last_event, tpd_I6_O, TRUE),
                 7 => (I7_ipd'last_event, tpd_I7_O, TRUE),
                 8 => (I8_ipd'last_event, tpd_I8_O, TRUE),
                 9 => (I9_ipd'last_event, tpd_I9_O, TRUE),
                 10 => (I10_ipd'last_event, tpd_I10_O, TRUE),
                 11 => (I11_ipd'last_event, tpd_I11_O, TRUE),
                 12 => (I12_ipd'last_event, tpd_I12_O, TRUE),
                 13 => (I13_ipd'last_event, tpd_I13_O, TRUE),
                 14 => (I14_ipd'last_event, tpd_I14_O, TRUE),
                 15 => (I15_ipd'last_event, tpd_I15_O, TRUE),
                 16 => (I16_ipd'last_event, tpd_I16_O, TRUE),
                 17 => (I17_ipd'last_event, tpd_I17_O, TRUE),
                 18 => (I18_ipd'last_event, tpd_I18_O, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;
 
configuration CFG_AND19_VITAL of AND19 is 
        for VITAL_VF
        end for; 
end CFG_AND19_VITAL;
----- VITAL model for cell AND2 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AND2 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_I0_O                       :	VitalDelayType01 := (1.25 ns, 1.25 ns);
      tpd_I1_O                       :	VitalDelayType01 := (1.25 ns, 1.25 ns);
      tipd_I0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      I0                             :	in    STD_ULOGIC;
      I1                             :	in    STD_ULOGIC;
      O                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AND2 : entity is TRUE;
end AND2;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library VF1;
architecture VITAL_VF of AND2 is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL I0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I1_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (I0_ipd, I0, tipd_I0);
   VitalWireDelay (I1_ipd, I1, tipd_I1);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (I0_ipd, I1_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS O_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE O_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      O_zd := (I1_ipd) AND (I0_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => O,
       GlitchData => O_GlitchData,
       OutSignalName => "O",
       OutTemp => O_zd,
       Paths => (0 => (I0_ipd'last_event, tpd_I0_O, TRUE),
                 1 => (I1_ipd'last_event, tpd_I1_O, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;

configuration CFG_AND2_VITAL of AND2 is 
        for VITAL_VF
        end for; 
end CFG_AND2_VITAL;
----- VITAL model for cell AND20 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AND20 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_I0_O                       :	VitalDelayType01 := (4.300 ns, 4.300 ns);
      tpd_I1_O                       :	VitalDelayType01 := (4.300 ns, 4.300 ns);
      tpd_I2_O                       :	VitalDelayType01 := (4.300 ns, 4.300 ns);
      tpd_I3_O                       :	VitalDelayType01 := (4.300 ns, 4.300 ns);
      tpd_I4_O                       :	VitalDelayType01 := (4.300 ns, 4.300 ns);
      tpd_I5_O                       :	VitalDelayType01 := (4.300 ns, 4.300 ns);
      tpd_I6_O                       :	VitalDelayType01 := (4.300 ns, 4.300 ns);
      tpd_I7_O                       :	VitalDelayType01 := (4.300 ns, 4.300 ns);
      tpd_I8_O                       :	VitalDelayType01 := (4.300 ns, 4.300 ns);
      tpd_I9_O                       :	VitalDelayType01 := (4.300 ns, 4.300 ns);
      tpd_I10_O                      :	VitalDelayType01 := (4.300 ns, 4.300 ns);
      tpd_I11_O                      :	VitalDelayType01 := (4.300 ns, 4.300 ns);
      tpd_I12_O                      :	VitalDelayType01 := (4.300 ns, 4.300 ns);
      tpd_I13_O                      :	VitalDelayType01 := (4.300 ns, 4.300 ns);
      tpd_I14_O                      :	VitalDelayType01 := (4.300 ns, 4.300 ns);
      tpd_I15_O                      :	VitalDelayType01 := (4.300 ns, 4.300 ns);
      tpd_I16_O                      :	VitalDelayType01 := (4.300 ns, 4.300 ns);
      tpd_I17_O                      :	VitalDelayType01 := (4.300 ns, 4.300 ns);
      tpd_I18_O                      :	VitalDelayType01 := (4.300 ns, 4.300 ns);
      tpd_I19_O                      :	VitalDelayType01 := (4.300 ns, 4.300 ns);
      tipd_I0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I2                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I3                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I4                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I5                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I6                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I7                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I8                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I9                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I10                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I11                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I12                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I13                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I14                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I15                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I16                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I17                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I18                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I19                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      I0                             :	in    STD_ULOGIC;
      I1                             :	in    STD_ULOGIC;
      I2                             :	in    STD_ULOGIC;
      I3                             :	in    STD_ULOGIC;
      I4                             :	in    STD_ULOGIC;
      I5                             :	in    STD_ULOGIC;
      I6                             :	in    STD_ULOGIC;
      I7                             :	in    STD_ULOGIC;
      I8                             :	in    STD_ULOGIC;
      I9                             :	in    STD_ULOGIC;
      I10                            :	in    STD_ULOGIC;
      I11                            :	in    STD_ULOGIC;
      I12                            :	in    STD_ULOGIC;
      I13                            :	in    STD_ULOGIC;
      I14                            :	in    STD_ULOGIC;
      I15                            :	in    STD_ULOGIC;
      I16                            :	in    STD_ULOGIC;
      I17                            :	in    STD_ULOGIC;
      I18                            :	in    STD_ULOGIC;
      I19                            :	in    STD_ULOGIC;
      O                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AND20 : entity is TRUE;
end AND20;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
 
library VF1;
architecture VITAL_VF of AND20 is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL I0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I1_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I2_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I3_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I4_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I5_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I6_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I7_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I8_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I9_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I10_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I11_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I12_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I13_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I14_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I15_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I16_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I17_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I18_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I19_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (I0_ipd, I0, tipd_I0);
   VitalWireDelay (I1_ipd, I1, tipd_I1);
   VitalWireDelay (I2_ipd, I2, tipd_I2);
   VitalWireDelay (I3_ipd, I3, tipd_I3);
   VitalWireDelay (I4_ipd, I4, tipd_I4);
   VitalWireDelay (I5_ipd, I5, tipd_I5);
   VitalWireDelay (I6_ipd, I6, tipd_I6);
   VitalWireDelay (I7_ipd, I7, tipd_I7);
   VitalWireDelay (I8_ipd, I8, tipd_I8);
   VitalWireDelay (I9_ipd, I9, tipd_I9);
   VitalWireDelay (I10_ipd, I10, tipd_I10);
   VitalWireDelay (I11_ipd, I11, tipd_I11);
   VitalWireDelay (I12_ipd, I12, tipd_I12);
   VitalWireDelay (I13_ipd, I13, tipd_I13);
   VitalWireDelay (I14_ipd, I14, tipd_I14);
   VitalWireDelay (I15_ipd, I15, tipd_I15);
   VitalWireDelay (I16_ipd, I16, tipd_I16);
   VitalWireDelay (I17_ipd, I17, tipd_I17);
   VitalWireDelay (I18_ipd, I18, tipd_I18);
   VitalWireDelay (I19_ipd, I19, tipd_I19);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (I0_ipd, I1_ipd, I2_ipd, I3_ipd, I4_ipd, I5_ipd, I6_ipd, I7_ipd, I8_ipd, I9_ipd, I10_ipd, I11_ipd, I12_ipd, I13_ipd, I14_ipd, I15_ipd, I16_ipd, I17_ipd, I18_ipd, I19_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS O_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE O_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      O_zd :=
       (I1_ipd) AND (I0_ipd) AND (I2_ipd) AND (I3_ipd) AND (I4_ipd) AND
         (I5_ipd) AND (I6_ipd) AND (I7_ipd) AND (I8_ipd) AND (I9_ipd) AND
         (I10_ipd) AND (I11_ipd) AND (I12_ipd) AND (I13_ipd) AND (I14_ipd)
         AND (I15_ipd) AND (I16_ipd) AND (I17_ipd) AND (I18_ipd) AND
         (I19_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => O,
       GlitchData => O_GlitchData,
       OutSignalName => "O",
       OutTemp => O_zd,
       Paths => (0 => (I0_ipd'last_event, tpd_I0_O, TRUE),
                 1 => (I1_ipd'last_event, tpd_I1_O, TRUE),
                 2 => (I2_ipd'last_event, tpd_I2_O, TRUE),
                 3 => (I3_ipd'last_event, tpd_I3_O, TRUE),
                 4 => (I4_ipd'last_event, tpd_I4_O, TRUE),
                 5 => (I5_ipd'last_event, tpd_I5_O, TRUE),
                 6 => (I6_ipd'last_event, tpd_I6_O, TRUE),
                 7 => (I7_ipd'last_event, tpd_I7_O, TRUE),
                 8 => (I8_ipd'last_event, tpd_I8_O, TRUE),
                 9 => (I9_ipd'last_event, tpd_I9_O, TRUE),
                 10 => (I10_ipd'last_event, tpd_I10_O, TRUE),
                 11 => (I11_ipd'last_event, tpd_I11_O, TRUE),
                 12 => (I12_ipd'last_event, tpd_I12_O, TRUE),
                 13 => (I13_ipd'last_event, tpd_I13_O, TRUE),
                 14 => (I14_ipd'last_event, tpd_I14_O, TRUE),
                 15 => (I15_ipd'last_event, tpd_I15_O, TRUE),
                 16 => (I16_ipd'last_event, tpd_I16_O, TRUE),
                 17 => (I17_ipd'last_event, tpd_I17_O, TRUE),
                 18 => (I18_ipd'last_event, tpd_I18_O, TRUE),
                 19 => (I19_ipd'last_event, tpd_I19_O, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;
 
configuration CFG_AND20_VITAL of AND20 is 
        for VITAL_VF
        end for; 
end CFG_AND20_VITAL;
----- VITAL model for cell AND3 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AND3 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_I0_O                       :	VitalDelayType01 := (1.25 ns, 1.25 ns);
      tpd_I1_O                       :	VitalDelayType01 := (1.25 ns, 1.25 ns);
      tpd_I2_O                       :	VitalDelayType01 := (1.25 ns, 1.25 ns);
      tipd_I0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I2                        :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      I0                             :	in    STD_ULOGIC;
      I1                             :	in    STD_ULOGIC;
      I2                             :	in    STD_ULOGIC;
      O                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AND3 : entity is TRUE;
end AND3;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library VF1;
architecture VITAL_VF of AND3 is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL I0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I1_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I2_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (I0_ipd, I0, tipd_I0);
   VitalWireDelay (I1_ipd, I1, tipd_I1);
   VitalWireDelay (I2_ipd, I2, tipd_I2);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (I0_ipd, I1_ipd, I2_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS O_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE O_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      O_zd := (I1_ipd) AND (I0_ipd) AND (I2_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => O,
       GlitchData => O_GlitchData,
       OutSignalName => "O",
       OutTemp => O_zd,
       Paths => (0 => (I0_ipd'last_event, tpd_I0_O, TRUE),
                 1 => (I1_ipd'last_event, tpd_I1_O, TRUE),
                 2 => (I2_ipd'last_event, tpd_I2_O, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;

configuration CFG_AND3_VITAL of AND3 is 
        for VITAL_VF
        end for; 
end CFG_AND3_VITAL;
----- VITAL model for cell AND4 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AND4 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_I0_O                       :	VitalDelayType01 := (1.80 ns, 1.80 ns);
      tpd_I1_O                       :	VitalDelayType01 := (1.80 ns, 1.80 ns);
      tpd_I2_O                       :	VitalDelayType01 := (1.80 ns, 1.80 ns);
      tpd_I3_O                       :	VitalDelayType01 := (1.80 ns, 1.80 ns);
      tipd_I0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I2                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I3                        :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      I0                             :	in    STD_ULOGIC;
      I1                             :	in    STD_ULOGIC;
      I2                             :	in    STD_ULOGIC;
      I3                             :	in    STD_ULOGIC;
      O                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AND4 : entity is TRUE;
end AND4;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library VF1;
architecture VITAL_VF of AND4 is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL I0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I1_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I2_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I3_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (I0_ipd, I0, tipd_I0);
   VitalWireDelay (I1_ipd, I1, tipd_I1);
   VitalWireDelay (I2_ipd, I2, tipd_I2);
   VitalWireDelay (I3_ipd, I3, tipd_I3);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (I0_ipd, I1_ipd, I2_ipd, I3_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS O_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE O_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      O_zd := (I1_ipd) AND (I0_ipd) AND (I2_ipd) AND (I3_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => O,
       GlitchData => O_GlitchData,
       OutSignalName => "O",
       OutTemp => O_zd,
       Paths => (0 => (I0_ipd'last_event, tpd_I0_O, TRUE),
                 1 => (I1_ipd'last_event, tpd_I1_O, TRUE),
                 2 => (I2_ipd'last_event, tpd_I2_O, TRUE),
                 3 => (I3_ipd'last_event, tpd_I3_O, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;

configuration CFG_AND4_VITAL of AND4 is 
        for VITAL_VF
        end for; 
end CFG_AND4_VITAL;
----- VITAL model for cell AND5 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AND5 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_I0_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I1_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I2_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I3_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I4_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tipd_I0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I2                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I3                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I4                        :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      I0                             :	in    STD_ULOGIC;
      I1                             :	in    STD_ULOGIC;
      I2                             :	in    STD_ULOGIC;
      I3                             :	in    STD_ULOGIC;
      I4                             :	in    STD_ULOGIC;
      O                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AND5 : entity is TRUE;
end AND5;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
 
library VF1;
architecture VITAL_VF of AND5 is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL I0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I1_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I2_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I3_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I4_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (I0_ipd, I0, tipd_I0);
   VitalWireDelay (I1_ipd, I1, tipd_I1);
   VitalWireDelay (I2_ipd, I2, tipd_I2);
   VitalWireDelay (I3_ipd, I3, tipd_I3);
   VitalWireDelay (I4_ipd, I4, tipd_I4);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (I0_ipd, I1_ipd, I2_ipd, I3_ipd, I4_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS O_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE O_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      O_zd :=
       (I1_ipd) AND (I0_ipd) AND (I2_ipd) AND (I3_ipd) AND (I4_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => O,
       GlitchData => O_GlitchData,
       OutSignalName => "O",
       OutTemp => O_zd,
       Paths => (0 => (I0_ipd'last_event, tpd_I0_O, TRUE),
                 1 => (I1_ipd'last_event, tpd_I1_O, TRUE),
                 2 => (I2_ipd'last_event, tpd_I2_O, TRUE),
                 3 => (I3_ipd'last_event, tpd_I3_O, TRUE),
                 4 => (I4_ipd'last_event, tpd_I4_O, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;
 
configuration CFG_AND5_VITAL of AND5 is 
        for VITAL_VF
        end for; 
end CFG_AND5_VITAL;
----- VITAL model for cell AND6 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AND6 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_I0_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I1_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I2_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I3_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I4_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I5_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tipd_I0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I2                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I3                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I4                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I5                        :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      I0                             :	in    STD_ULOGIC;
      I1                             :	in    STD_ULOGIC;
      I2                             :	in    STD_ULOGIC;
      I3                             :	in    STD_ULOGIC;
      I4                             :	in    STD_ULOGIC;
      I5                             :	in    STD_ULOGIC;
      O                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AND6 : entity is TRUE;
end AND6;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
 
library VF1;
architecture VITAL_VF of AND6 is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL I0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I1_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I2_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I3_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I4_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I5_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (I0_ipd, I0, tipd_I0);
   VitalWireDelay (I1_ipd, I1, tipd_I1);
   VitalWireDelay (I2_ipd, I2, tipd_I2);
   VitalWireDelay (I3_ipd, I3, tipd_I3);
   VitalWireDelay (I4_ipd, I4, tipd_I4);
   VitalWireDelay (I5_ipd, I5, tipd_I5);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (I0_ipd, I1_ipd, I2_ipd, I3_ipd, I4_ipd, I5_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS O_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE O_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      O_zd :=
       (I1_ipd) AND (I0_ipd) AND (I2_ipd) AND (I3_ipd) AND (I4_ipd) AND
         (I5_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => O,
       GlitchData => O_GlitchData,
       OutSignalName => "O",
       OutTemp => O_zd,
       Paths => (0 => (I0_ipd'last_event, tpd_I0_O, TRUE),
                 1 => (I1_ipd'last_event, tpd_I1_O, TRUE),
                 2 => (I2_ipd'last_event, tpd_I2_O, TRUE),
                 3 => (I3_ipd'last_event, tpd_I3_O, TRUE),
                 4 => (I4_ipd'last_event, tpd_I4_O, TRUE),
                 5 => (I5_ipd'last_event, tpd_I5_O, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;
 
configuration CFG_AND6_VITAL of AND6 is 
        for VITAL_VF
        end for; 
end CFG_AND6_VITAL;
----- VITAL model for cell AND7 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AND7 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_I0_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I1_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I2_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I3_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I4_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I5_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I6_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tipd_I0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I2                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I3                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I4                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I5                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I6                        :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      I0                             :	in    STD_ULOGIC;
      I1                             :	in    STD_ULOGIC;
      I2                             :	in    STD_ULOGIC;
      I3                             :	in    STD_ULOGIC;
      I4                             :	in    STD_ULOGIC;
      I5                             :	in    STD_ULOGIC;
      I6                             :	in    STD_ULOGIC;
      O                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AND7 : entity is TRUE;
end AND7;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
 
library VF1;
architecture VITAL_VF of AND7 is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL I0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I1_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I2_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I3_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I4_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I5_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I6_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (I0_ipd, I0, tipd_I0);
   VitalWireDelay (I1_ipd, I1, tipd_I1);
   VitalWireDelay (I2_ipd, I2, tipd_I2);
   VitalWireDelay (I3_ipd, I3, tipd_I3);
   VitalWireDelay (I4_ipd, I4, tipd_I4);
   VitalWireDelay (I5_ipd, I5, tipd_I5);
   VitalWireDelay (I6_ipd, I6, tipd_I6);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (I0_ipd, I1_ipd, I2_ipd, I3_ipd, I4_ipd, I5_ipd, I6_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS O_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE O_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      O_zd :=
       (I1_ipd) AND (I0_ipd) AND (I2_ipd) AND (I3_ipd) AND (I4_ipd) AND
         (I5_ipd) AND (I6_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => O,
       GlitchData => O_GlitchData,
       OutSignalName => "O",
       OutTemp => O_zd,
       Paths => (0 => (I0_ipd'last_event, tpd_I0_O, TRUE),
                 1 => (I1_ipd'last_event, tpd_I1_O, TRUE),
                 2 => (I2_ipd'last_event, tpd_I2_O, TRUE),
                 3 => (I3_ipd'last_event, tpd_I3_O, TRUE),
                 4 => (I4_ipd'last_event, tpd_I4_O, TRUE),
                 5 => (I5_ipd'last_event, tpd_I5_O, TRUE),
                 6 => (I6_ipd'last_event, tpd_I6_O, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;
 
configuration CFG_AND7_VITAL of AND7 is 
        for VITAL_VF
        end for; 
end CFG_AND7_VITAL;
----- VITAL model for cell AND8 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AND8 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_I0_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I1_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I2_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I3_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I4_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I5_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I6_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I7_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tipd_I0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I2                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I3                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I4                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I5                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I6                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I7                        :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      I0                             :	in    STD_ULOGIC;
      I1                             :	in    STD_ULOGIC;
      I2                             :	in    STD_ULOGIC;
      I3                             :	in    STD_ULOGIC;
      I4                             :	in    STD_ULOGIC;
      I5                             :	in    STD_ULOGIC;
      I6                             :	in    STD_ULOGIC;
      I7                             :	in    STD_ULOGIC;
      O                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AND8 : entity is TRUE;
end AND8;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
 
library VF1;
architecture VITAL_VF of AND8 is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL I0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I1_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I2_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I3_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I4_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I5_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I6_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I7_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (I0_ipd, I0, tipd_I0);
   VitalWireDelay (I1_ipd, I1, tipd_I1);
   VitalWireDelay (I2_ipd, I2, tipd_I2);
   VitalWireDelay (I3_ipd, I3, tipd_I3);
   VitalWireDelay (I4_ipd, I4, tipd_I4);
   VitalWireDelay (I5_ipd, I5, tipd_I5);
   VitalWireDelay (I6_ipd, I6, tipd_I6);
   VitalWireDelay (I7_ipd, I7, tipd_I7);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (I0_ipd, I1_ipd, I2_ipd, I3_ipd, I4_ipd, I5_ipd, I6_ipd, I7_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS O_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE O_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      O_zd :=
       (I1_ipd) AND (I0_ipd) AND (I2_ipd) AND (I3_ipd) AND (I4_ipd) AND
         (I5_ipd) AND (I6_ipd) AND (I7_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => O,
       GlitchData => O_GlitchData,
       OutSignalName => "O",
       OutTemp => O_zd,
       Paths => (0 => (I0_ipd'last_event, tpd_I0_O, TRUE),
                 1 => (I1_ipd'last_event, tpd_I1_O, TRUE),
                 2 => (I2_ipd'last_event, tpd_I2_O, TRUE),
                 3 => (I3_ipd'last_event, tpd_I3_O, TRUE),
                 4 => (I4_ipd'last_event, tpd_I4_O, TRUE),
                 5 => (I5_ipd'last_event, tpd_I5_O, TRUE),
                 6 => (I6_ipd'last_event, tpd_I6_O, TRUE),
                 7 => (I7_ipd'last_event, tpd_I7_O, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;
 
configuration CFG_AND8_VITAL of AND8 is 
        for VITAL_VF
        end for; 
end CFG_AND8_VITAL;
----- VITAL model for cell AND9 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AND9 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_I0_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I1_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I2_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I3_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I4_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I5_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I6_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I7_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I8_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tipd_I0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I2                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I3                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I4                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I5                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I6                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I7                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I8                        :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      I0                             :	in    STD_ULOGIC;
      I1                             :	in    STD_ULOGIC;
      I2                             :	in    STD_ULOGIC;
      I3                             :	in    STD_ULOGIC;
      I4                             :	in    STD_ULOGIC;
      I5                             :	in    STD_ULOGIC;
      I6                             :	in    STD_ULOGIC;
      I7                             :	in    STD_ULOGIC;
      I8                             :	in    STD_ULOGIC;
      O                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AND9 : entity is TRUE;
end AND9;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
 
library VF1;
architecture VITAL_VF of AND9 is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL I0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I1_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I2_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I3_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I4_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I5_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I6_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I7_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I8_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (I0_ipd, I0, tipd_I0);
   VitalWireDelay (I1_ipd, I1, tipd_I1);
   VitalWireDelay (I2_ipd, I2, tipd_I2);
   VitalWireDelay (I3_ipd, I3, tipd_I3);
   VitalWireDelay (I4_ipd, I4, tipd_I4);
   VitalWireDelay (I5_ipd, I5, tipd_I5);
   VitalWireDelay (I6_ipd, I6, tipd_I6);
   VitalWireDelay (I7_ipd, I7, tipd_I7);
   VitalWireDelay (I8_ipd, I8, tipd_I8);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (I0_ipd, I1_ipd, I2_ipd, I3_ipd, I4_ipd, I5_ipd, I6_ipd, I7_ipd, I8_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS O_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE O_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      O_zd :=
       (I1_ipd) AND (I0_ipd) AND (I2_ipd) AND (I3_ipd) AND (I4_ipd) AND
         (I5_ipd) AND (I6_ipd) AND (I7_ipd) AND (I8_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => O,
       GlitchData => O_GlitchData,
       OutSignalName => "O",
       OutTemp => O_zd,
       Paths => (0 => (I0_ipd'last_event, tpd_I0_O, TRUE),
                 1 => (I1_ipd'last_event, tpd_I1_O, TRUE),
                 2 => (I2_ipd'last_event, tpd_I2_O, TRUE),
                 3 => (I3_ipd'last_event, tpd_I3_O, TRUE),
                 4 => (I4_ipd'last_event, tpd_I4_O, TRUE),
                 5 => (I5_ipd'last_event, tpd_I5_O, TRUE),
                 6 => (I6_ipd'last_event, tpd_I6_O, TRUE),
                 7 => (I7_ipd'last_event, tpd_I7_O, TRUE),
                 8 => (I8_ipd'last_event, tpd_I8_O, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;
 
configuration CFG_AND9_VITAL of AND9 is 
        for VITAL_VF
        end for; 
end CFG_AND9_VITAL;
----- VITAL model for cell AO21 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AO21 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_I0_O                       :	VitalDelayType01 := (1.25 ns, 1.25 ns);
      tpd_I1_O                       :	VitalDelayType01 := (1.25 ns, 1.25 ns);
      tpd_I2_O                       :	VitalDelayType01 := (1.25 ns, 1.25 ns);
      tipd_I0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I2                        :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      I0                             :	in    STD_ULOGIC;
      I1                             :	in    STD_ULOGIC;
      I2                             :	in    STD_ULOGIC;
      O                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AO21 : entity is TRUE;
end AO21;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library VF1;
architecture VITAL_VF of AO21 is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL I0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I1_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I2_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (I0_ipd, I0, tipd_I0);
   VitalWireDelay (I1_ipd, I1, tipd_I1);
   VitalWireDelay (I2_ipd, I2, tipd_I2);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (I0_ipd, I1_ipd, I2_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS O_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE O_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      O_zd := (I2_ipd) OR ((I1_ipd) AND (I0_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => O,
       GlitchData => O_GlitchData,
       OutSignalName => "O",
       OutTemp => O_zd,
       Paths => (0 => (I0_ipd'last_event, tpd_I0_O, TRUE),
                 1 => (I1_ipd'last_event, tpd_I1_O, TRUE),
                 2 => (I2_ipd'last_event, tpd_I2_O, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;

configuration CFG_AO21_VITAL of AO21 is 
        for VITAL_VF
        end for; 
end CFG_AO21_VITAL;
----- VITAL model for cell AO221 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AO221 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_I0_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I1_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I2_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I3_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I4_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tipd_I0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I2                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I3                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I4                        :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      I0                             :	in    STD_ULOGIC;
      I1                             :	in    STD_ULOGIC;
      I2                             :	in    STD_ULOGIC;
      I3                             :	in    STD_ULOGIC;
      I4                             :	in    STD_ULOGIC;
      O                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AO221 : entity is TRUE;
end AO221;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
 
library VF1;
architecture VITAL_VF of AO221 is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL I0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I1_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I2_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I3_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I4_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (I0_ipd, I0, tipd_I0);
   VitalWireDelay (I1_ipd, I1, tipd_I1);
   VitalWireDelay (I2_ipd, I2, tipd_I2);
   VitalWireDelay (I3_ipd, I3, tipd_I3);
   VitalWireDelay (I4_ipd, I4, tipd_I4);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (I0_ipd, I1_ipd, I2_ipd, I3_ipd, I4_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS O_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE O_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      O_zd :=
       ((I3_ipd) AND (I2_ipd)) OR ((I1_ipd) AND (I0_ipd)) OR (I4_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => O,
       GlitchData => O_GlitchData,
       OutSignalName => "O",
       OutTemp => O_zd,
       Paths => (0 => (I0_ipd'last_event, tpd_I0_O, TRUE),
                 1 => (I1_ipd'last_event, tpd_I1_O, TRUE),
                 2 => (I2_ipd'last_event, tpd_I2_O, TRUE),
                 3 => (I3_ipd'last_event, tpd_I3_O, TRUE),
                 4 => (I4_ipd'last_event, tpd_I4_O, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;
 
configuration CFG_AO221_VITAL of AO221 is 
        for VITAL_VF
        end for; 
end CFG_AO221_VITAL;
----- VITAL model for cell AO321 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AO321 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_I0_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I1_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I2_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I3_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I4_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I5_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tipd_I0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I2                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I3                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I4                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I5                        :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      I0                             :	in    STD_ULOGIC;
      I1                             :	in    STD_ULOGIC;
      I2                             :	in    STD_ULOGIC;
      I3                             :	in    STD_ULOGIC;
      I4                             :	in    STD_ULOGIC;
      I5                             :	in    STD_ULOGIC;
      O                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AO321 : entity is TRUE;
end AO321;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library VF1;
architecture VITAL_VF of AO321 is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL I0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I1_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I2_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I3_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I4_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I5_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (I0_ipd, I0, tipd_I0);
   VitalWireDelay (I1_ipd, I1, tipd_I1);
   VitalWireDelay (I2_ipd, I2, tipd_I2);
   VitalWireDelay (I3_ipd, I3, tipd_I3);
   VitalWireDelay (I4_ipd, I4, tipd_I4);
   VitalWireDelay (I5_ipd, I5, tipd_I5);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (I0_ipd, I1_ipd, I2_ipd, I3_ipd, I4_ipd, I5_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS O_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE O_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      O_zd :=
       ((I4_ipd) AND (I3_ipd)) OR ((I1_ipd) AND (I0_ipd) AND (I2_ipd)) OR
         (I5_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => O,
       GlitchData => O_GlitchData,
       OutSignalName => "O",
       OutTemp => O_zd,
       Paths => (0 => (I0_ipd'last_event, tpd_I0_O, TRUE),
                 1 => (I1_ipd'last_event, tpd_I1_O, TRUE),
                 2 => (I2_ipd'last_event, tpd_I2_O, TRUE),
                 3 => (I3_ipd'last_event, tpd_I3_O, TRUE),
                 4 => (I4_ipd'last_event, tpd_I4_O, TRUE),
                 5 => (I5_ipd'last_event, tpd_I5_O, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;

configuration CFG_AO321_VITAL of AO321 is 
        for VITAL_VF
        end for; 
end CFG_AO321_VITAL;
----- VITAL model for cell AS_LSB -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AS_LSB is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_A0_S0                      :	VitalDelayType01 := (1.800 ns, 1.800 ns);
      tpd_B0_S0                      :	VitalDelayType01 := (1.800 ns, 1.800 ns);
      tpd_CIN_S0                     :	VitalDelayType01 := (1.800 ns, 1.800 ns);
      tpd_AS_S0                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A0_COUT                    :	VitalDelayType01 := (1.800 ns, 1.800 ns);
      tpd_B0_COUT                    :	VitalDelayType01 := (1.800 ns, 1.800 ns);
      tpd_CIN_COUT                   :	VitalDelayType01 := (0.200 ns, 0.200 ns);
      tpd_AS_COUT                    :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CIN                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_AS                        :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A0                             :	in    STD_ULOGIC;
      B0                             :	in    STD_ULOGIC;
      CIN                            :	in    STD_ULOGIC;
      AS                             :	in    STD_ULOGIC;
      S0                             :	out   STD_ULOGIC;
      COUT                           :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AS_LSB : entity is TRUE;
end AS_LSB;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library VF1;
architecture VITAL_VF of AS_LSB is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL A0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CIN_ipd	 : STD_ULOGIC := 'X';
   SIGNAL AS_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A0_ipd, A0, tipd_A0);
   VitalWireDelay (B0_ipd, B0, tipd_B0);
   VitalWireDelay (CIN_ipd, CIN, tipd_CIN);
   VitalWireDelay (AS_ipd, AS, tipd_AS);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A0_ipd, B0_ipd, CIN_ipd, AS_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS S0_zd : STD_LOGIC is Results(1);
   ALIAS COUT_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE S0_GlitchData	: VitalGlitchDataType;
   VARIABLE COUT_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      S0_zd := (B0_ipd) XOR (A0_ipd) XOR (CIN_ipd);
      COUT_zd :=
       (((NOT ((AS_ipd) XOR (CIN_ipd)))) AND (A0_ipd)) OR (((NOT ((AS_ipd)
         XOR (B0_ipd)))) AND (A0_ipd)) OR (((NOT ((AS_ipd) XOR (CIN_ipd))))
         AND ((NOT ((AS_ipd) XOR (B0_ipd)))));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => S0,
       GlitchData => S0_GlitchData,
       OutSignalName => "S0",
       OutTemp => S0_zd,
       Paths => (0 => (A0_ipd'last_event, tpd_A0_S0, TRUE),
                 1 => (B0_ipd'last_event, tpd_B0_S0, TRUE),
                 2 => (CIN_ipd'last_event, tpd_CIN_S0, TRUE),
                 3 => (AS_ipd'last_event, tpd_AS_S0, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);
      VitalPathDelay01 (
       OutSignal => COUT,
       GlitchData => COUT_GlitchData,
       OutSignalName => "COUT",
       OutTemp => COUT_zd,
       Paths => (0 => (A0_ipd'last_event, tpd_A0_COUT, TRUE),
                 1 => (B0_ipd'last_event, tpd_B0_COUT, TRUE),
                 2 => (CIN_ipd'last_event, tpd_CIN_COUT, TRUE),
                 3 => (AS_ipd'last_event, tpd_AS_COUT, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;

configuration CFG_AS_LSB_VITAL of AS_LSB is 
        for VITAL_VF
        end for; 
end CFG_AS_LSB_VITAL;
----- VITAL model for cell BIPAD -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


----- VITAL model for cell BI_DIR -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity BI_DIR is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_OE_IO                      :	VitalDelayType01Z := (0.640 ns, 0.640 ns, 0.640 ns, 0.640 ns, 0.640 ns, 0.640 ns);
      tpd_I0_IO                      :	VitalDelayType01 := (0.640 ns, 0.640 ns);
      tpd_IO_O                       :	VitalDelayType01 := (0.400 ns, 0.400 ns);
      tipd_I0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_OE                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_IO                        :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      I0                             :	in    STD_ULOGIC;
      OE                             :	in    STD_ULOGIC;
      IO                             :	inout STD_ULOGIC;
      O                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of BI_DIR : entity is TRUE;
end BI_DIR;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library VF1;
--use VF1.VTABLES.all;
architecture VITAL_VF of BI_DIR is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL I0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL OE_ipd	 : STD_ULOGIC := 'X';
   SIGNAL IO_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (I0_ipd, I0, tipd_I0);
   VitalWireDelay (OE_ipd, OE, tipd_OE);
   VitalWireDelay (IO_ipd, IO, tipd_IO);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (I0_ipd, OE_ipd, IO_ipd)


   -- functionality results
--   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
     VARIABLE IO_zd : std_ulogic ;
     VARIABLE O_zd : std_ulogic ;

   -- output glitch detection variables
   VARIABLE IO_GlitchData	: VitalGlitchDataType;
   VARIABLE O_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      IO_zd := VitalBUFIF1 (I0_ipd, OE_ipd);
      O_zd := VitalBUF(IO_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01Z (
       OutSignal => IO,
       GlitchData => IO_GlitchData,
       OutSignalName => "IO",
       OutTemp => IO_zd,
       Paths => (0 => (OE_ipd'last_event, VitalExtendToFillDelay(tpd_OE_IO), TRUE),
                 1 => (I0_ipd'last_event, VitalExtendToFillDelay(tpd_I0_IO), TRUE)),
       Mode => VitalInertial,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING,
       OutputMap => "UX01ZWLH-");
      VitalPathDelay01 (
       OutSignal => O,
       GlitchData => O_GlitchData,
       OutSignalName => "O",
       OutTemp => O_zd,
       Paths => (0 => (IO_ipd'last_event, tpd_IO_O, TRUE)),
       Mode => VitalInertial,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;

configuration CFG_BI_DIR_VITAL of BI_DIR is 
        for VITAL_VF
        end for; 
end CFG_BI_DIR_VITAL;
----- VITAL model for cell BUFF -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity BUFF is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_I0_O                       :	VitalDelayType01 := (1.25 ns, 1.25 ns);
      tipd_I0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      I0                             :	in    STD_ULOGIC;
      O                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of BUFF : entity is TRUE;
end BUFF;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library VF1;
architecture VITAL_VF of BUFF is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL I0_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (I0_ipd, I0, tipd_I0);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (I0_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS O_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE O_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      O_zd := TO_X01(I0_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => O,
       GlitchData => O_GlitchData,
       OutSignalName => "O",
       OutTemp => O_zd,
       Paths => (0 => (I0_ipd'last_event, tpd_I0_O, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;

configuration CFG_BUFF_VITAL of BUFF is 
        for VITAL_VF
        end for; 
end CFG_BUFF_VITAL;
----- VITAL model for cell BUFTH -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity BUFTH is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_OE_O                       :	VitalDelayType01Z := (0.640 ns, 0.640 ns, 0.640 ns, 0.640 ns, 0.640 ns, 0.640 ns);
      tpd_I0_O                       :	VitalDelayType01 := (0.640 ns, 0.640 ns);
      tipd_I0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_OE                        :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      I0                             :	in    STD_ULOGIC;
      OE                             :	in    STD_ULOGIC;
      O                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of BUFTH : entity is TRUE;
end BUFTH;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library VF1;
--use VF1.VTABLES.all;
architecture VITAL_VF of BUFTH is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL I0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL OE_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (I0_ipd, I0, tipd_I0);
   VitalWireDelay (OE_ipd, OE, tipd_OE);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (I0_ipd, OE_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS O_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE O_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      O_zd := VitalBUFIF0 (data => I0_ipd,
              enable => (NOT OE_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01Z (
       OutSignal => O,
       GlitchData => O_GlitchData,
       OutSignalName => "O",
       OutTemp => O_zd,
       Paths => (0 => (OE_ipd'last_event, VitalExtendToFillDelay(tpd_OE_O), TRUE),
                 1 => (I0_ipd'last_event, VitalExtendToFillDelay(tpd_I0_O), TRUE)),
       Mode => VitalInertial,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING,
       OutputMap => "UX01ZWLH-");

end process;
end VITAL_VF;

configuration CFG_BUFTH_VITAL of BUFTH is 
        for VITAL_VF
        end for; 
end CFG_BUFTH_VITAL;
----- VITAL model for cell BUFTI -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;
LIBRARY VF1 ;
use VF1.VLOGTOVITAL_TABLES.all;

-- entity declaration --
entity BUFTI is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_OE_O                       :	VitalDelayType01z := 
               (0.640 ns, 0.640 ns, 0.640 ns, 0.640 ns, 0.640 ns, 0.640 ns);
      tpd_I0_O                       :	VitalDelayType01 := (0.640 ns, 0.640 ns);
      tipd_I0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_OE                        :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      I0                             :	in    STD_ULOGIC;
      OE                             :	in    STD_ULOGIC;
      O                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of BUFTI : entity is TRUE;
end BUFTI;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library VF1;
architecture VITAL_VF of BUFTI is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL I0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL OE_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (I0_ipd, I0, tipd_I0);
   VitalWireDelay (OE_ipd, OE, tipd_OE);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (I0_ipd, OE_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS O_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE O_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      O_zd := VitalBUFIF0 (data => I0_ipd,
              enable => (NOT OE_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01Z (
       OutSignal => O,
       GlitchData => O_GlitchData,
       OutSignalName => "O",
       OutTemp => O_zd,
       Paths => (0 => (OE_ipd'last_event, VitalExtendToFillDelay(tpd_OE_O), TRUE),
                 1 => (I0_ipd'last_event, VitalExtendToFillDelay(tpd_I0_O), TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING,
       OutputMap => "UX01ZWLH-");

end process;
end VITAL_VF;

configuration CFG_BUFTI_VITAL of BUFTI is 
        for VITAL_VF
        end for; 
end CFG_BUFTI_VITAL;
----- VITAL model for cell BUFTL -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity BUFTL is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_OE_O                       :	VitalDelayType01Z := (0.640 ns, 0.640 ns, 0.640 ns, 0.640 ns, 0.640 ns, 0.640 ns);
      tpd_I0_O                       :	VitalDelayType01 := (0.640 ns, 0.640 ns);
      tipd_I0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_OE                        :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      I0                             :	in    STD_ULOGIC;
      OE                             :	in    STD_ULOGIC;
      O                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of BUFTL : entity is TRUE;
end BUFTL;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library VF1;
--use VF1.VTABLES.all;
architecture VITAL_VF of BUFTL is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL I0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL OE_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (I0_ipd, I0, tipd_I0);
   VitalWireDelay (OE_ipd, OE, tipd_OE);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (I0_ipd, OE_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS O_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE O_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      O_zd := VitalBUFIF0 (data => I0_ipd,
              enable => OE_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01Z (
       OutSignal => O,
       GlitchData => O_GlitchData,
       OutSignalName => "O",
       OutTemp => O_zd,
       Paths => (0 => (OE_ipd'last_event, VitalExtendToFillDelay(tpd_OE_O), TRUE),
                 1 => (I0_ipd'last_event, VitalExtendToFillDelay(tpd_I0_O), TRUE)),
       Mode => VitalInertial,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING,
       OutputMap => "UX01ZWLH-");

end process;
end VITAL_VF;

configuration CFG_BUFTL_VITAL of BUFTL is 
        for VITAL_VF
        end for; 
end CFG_BUFTL_VITAL;
---------------------------------------------------------------------------------
-- VITAL model for cell CCU_ABS
---------------------------------------------------------------------------------
LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.VITAL_timing.all;
USE IEEE.VITAL_primitives.all;
LIBRARY VF1;
USE VF1.all;
-----------------------------------------------------------------------------
--ENTITY DECLARATION
-----------------------------------------------------------------------------
ENTITY CCU_ABS IS

GENERIC (
	tipd_D			 : VITALDELAYTYPE01Z 	 := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
	tipd_PN			 : VITALDELAYTYPE01Z 	 := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
	tipd_CIN		 : VITALDELAYTYPE01Z 	 := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
	tpd_D_S0		 : VITALDELAYTYPE01 	 := (1.25 ns, 1.25 ns);
	tpd_PN_S0		 : VITALDELAYTYPE01 	 := (1.25 ns, 1.25 ns);
	tpd_CIN_S0		 : VITALDELAYTYPE01 	 := (1.25 ns, 1.25 ns);
	tpd_D_COUT		 : VITALDELAYTYPE01 	 := (1.25 ns, 1.25 ns);
	tpd_PN_COUT		 : VITALDELAYTYPE01 	 := (1.25 ns, 1.25 ns);
	tpd_CIN_COUT		 : VITALDELAYTYPE01 	 := (1.25 ns, 1.25 ns)
	);

PORT    (
	S0			 : OUT   std_logic;
	COUT			 : OUT   std_logic;
	D			 : IN    std_logic := 'U';
	PN			 : IN    std_logic := 'U';
	CIN			 : IN    std_logic := 'U'
	);

ATTRIBUTE VITAL_LEVEL0 OF CCU_ABS : ENTITY IS TRUE ;

END CCU_ABS;

-----------------------------------------------------------------------------
-- ARCHITECTURE declaration
-----------------------------------------------------------------------------
library IEEE;
use IEEE.VITAL_Primitives.all;
library VF1;
use VF1.all;
ARCHITECTURE VITAL_VF OF CCU_ABS  IS
	ATTRIBUTE VITAL_LEVEL1 OF VITAL_VF : ARCHITECTURE IS TRUE;

	SIGNAL	D_ipd			 : std_logic         := 'X';
	SIGNAL	PN_ipd			 : std_logic         := 'X';
	SIGNAL	CIN_ipd			 : std_logic         := 'X';
BEGIN
-----------------------------------------------------------------------------
-- INPUT PATH DELAYs
-----------------------------------------------------------------------------
WIREDELAY : BLOCK
BEGIN
	VitalWireDelay( D_ipd, D, tipd_D );
	VitalWireDelay( PN_ipd, PN, tipd_PN );
	VitalWireDelay( CIN_ipd, CIN, tipd_CIN );
END BLOCK;

-----------------------------------------------------------------------------
-- Behavior Section
-----------------------------------------------------------------------------

VitalBehaviour_0 : PROCESS(PN_ipd,D_ipd,CIN_ipd)

VARIABLE 	pn_zd			 : std_ulogic;
VARIABLE 	o1_zd			 : std_ulogic;
VARIABLE 	d_zd			 : std_ulogic;
VARIABLE 	cin_zd			 : std_ulogic;
VARIABLE 	o2_zd			 : std_ulogic;
VARIABLE 	S0_zd			 : std_ulogic;
VARIABLE 	o3_zd			 : std_ulogic;
VARIABLE 	COUT_zd			 : std_ulogic;
VARIABLE 	S0GLITCH_DATA		 : VitalGlitchDataType;
VARIABLE 	COUTGLITCH_DATA		 : VitalGlitchDataType;


BEGIN


--Functionality Section

pn_zd		 := VitalINV(PN_ipd);
o1_zd		 := VitalAND2(pn_zd,D_ipd);
d_zd		 := VitalINV(D_ipd);
cin_zd		 := VitalXOR2(d_zd,CIN_ipd);
o2_zd		 := VitalAND2(pn_ipd,cin_zd);
S0_zd		 := VitalOR2(o1_zd,o2_zd);
o3_zd		 := VitalAND2(d_zd,CIN_ipd);
COUT_zd		 := VitalAND2(PN_ipd,o3_zd);

--PathDelay Section

 VitalPathDelay01 ( S0, S0GLITCH_DATA, "S0", S0_zd,
	Paths => (
	0 => ( D_ipd'LAST_EVENT, tpd_D_S0, TRUE ),
	1 => ( PN_ipd'LAST_EVENT, tpd_PN_S0, TRUE ),
	2 => ( CIN_ipd'LAST_EVENT, tpd_CIN_S0, TRUE ) ),
	DefaultDelay=>VitalZeroDelay01,
	Mode=>VitalInertial,
	XON=>TRUE,
	MsgOn=>TRUE,
	MsgSeverity=>WARNING );

 VitalPathDelay01 ( COUT, COUTGLITCH_DATA, "COUT", COUT_zd,
	Paths => (
	0 => ( D_ipd'LAST_EVENT, tpd_D_COUT, TRUE ),
	1 => ( PN_ipd'LAST_EVENT, tpd_PN_COUT, TRUE ),
	2 => ( CIN_ipd'LAST_EVENT, tpd_CIN_COUT, TRUE ) ),
	DefaultDelay=>VitalZeroDelay01,
	Mode=>VitalInertial,
	XON=>TRUE,
	MsgOn=>TRUE,
	MsgSeverity=>WARNING );


END PROCESS VitalBehaviour_0;


END VITAL_VF;
configuration CFG_CCU_ABS_VITAL of CCU_ABS is 
        for VITAL_VF
        end for; 
end CFG_CCU_ABS_VITAL;
---------------------------------------------------------------------------------
-- VITAL model for cell CCU_AGB
---------------------------------------------------------------------------------
LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.VITAL_timing.all;
USE IEEE.VITAL_primitives.all;
LIBRARY VF1;
USE VF1.all;
-----------------------------------------------------------------------------
--ENTITY DECLARATION
-----------------------------------------------------------------------------
ENTITY CCU_AGB IS

GENERIC (
	tipd_A0			 : VITALDELAYTYPE01Z 	 := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
	tipd_B0			 : VITALDELAYTYPE01Z 	 := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
	tipd_CIN		 : VITALDELAYTYPE01Z 	 := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
	tpd_A0_COUT		 : VITALDELAYTYPE01 	 := (1.25 ns, 1.25 ns);
	tpd_B0_COUT		 : VITALDELAYTYPE01 	 := (1.25 ns, 1.25 ns);
	tpd_CIN_COUT		 : VITALDELAYTYPE01 	 := (1.25 ns, 1.25 ns)
	);

PORT    (
	COUT			 : OUT   std_logic;
	A0			 : IN    std_logic := 'U';
	B0			 : IN    std_logic := 'U';
	CIN			 : IN    std_logic := 'U'
	);

ATTRIBUTE VITAL_LEVEL0 OF CCU_AGB : ENTITY IS TRUE ;

END CCU_AGB;

-----------------------------------------------------------------------------
-- ARCHITECTURE declaration
-----------------------------------------------------------------------------
library IEEE;
use IEEE.VITAL_Primitives.all;
library VF1;
use VF1.all;
ARCHITECTURE VITAL_VF OF CCU_AGB  IS
	ATTRIBUTE VITAL_LEVEL1 OF VITAL_VF : ARCHITECTURE IS TRUE;

	SIGNAL	A0_ipd			 : std_logic         := 'X';
	SIGNAL	B0_ipd			 : std_logic         := 'X';
	SIGNAL	CIN_ipd			 : std_logic         := 'X';
BEGIN
-----------------------------------------------------------------------------
-- INPUT PATH DELAYs
-----------------------------------------------------------------------------
WIREDELAY : BLOCK
BEGIN
	VitalWireDelay( A0_ipd, A0, tipd_A0 );
	VitalWireDelay( B0_ipd, B0, tipd_B0 );
	VitalWireDelay( CIN_ipd, CIN, tipd_CIN );
END BLOCK;

-----------------------------------------------------------------------------
-- Behavior Section
-----------------------------------------------------------------------------

VitalBehaviour_0 : PROCESS(B0_ipd,A0_ipd,CIN_ipd)

VARIABLE 	b_zd			 : std_ulogic;
VARIABLE 	a_zd			 : std_ulogic;
VARIABLE 	a1_zd			 : std_ulogic;
VARIABLE 	a2_zd			 : std_ulogic;
VARIABLE 	COUT_zd			 : std_ulogic;
VARIABLE 	COUTGLITCH_DATA		 : VitalGlitchDataType;


BEGIN


--Functionality Section

b_zd		 := VitalINV(B0_ipd);
a_zd		 := VitalAND2(A0_ipd,b_zd);
a1_zd		 := VitalXNOR2(A0_ipd,B0_ipd);
a2_zd		 := VitalAND2(a1_zd,CIN_ipd);
COUT_zd		 := VitalOR2(a_zd,a2_zd);

--PathDelay Section

 VitalPathDelay01 (COUT,COUTGLITCH_DATA,"COUT",COUT_zd,
	Paths => (
	0 => ( A0_ipd'LAST_EVENT, tpd_A0_COUT, TRUE ),
	1 => ( B0_ipd'LAST_EVENT, tpd_B0_COUT, TRUE ),
	2 => ( CIN_ipd'LAST_EVENT, tpd_CIN_COUT, TRUE ) ),
	DefaultDelay=>VitalZeroDelay01,
	Mode=>VitalInertial,
	XON=>TRUE,
	MsgOn=>TRUE,
	MsgSeverity=>WARNING );


END PROCESS;
end VITAL_VF;
configuration CFG_CCU_AGB_VITAL of CCU_AGB is 
        for VITAL_VF
        end for; 
end CFG_CCU_AGB_VITAL;
---------------------------------------------------------------------------------
-- VITAL model for cell CCU_AS
---------------------------------------------------------------------------------
LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.VITAL_timing.all;
USE IEEE.VITAL_primitives.all;
LIBRARY VF1;
USE VF1.all;
-----------------------------------------------------------------------------
--ENTITY DECLARATION
-----------------------------------------------------------------------------
ENTITY CCU_AS IS

GENERIC (
	tipd_A0			 : VITALDELAYTYPE01Z 	 := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
	tipd_B0			 : VITALDELAYTYPE01Z 	 := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
	tipd_CIN		 : VITALDELAYTYPE01Z 	 := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
	tipd_AS			 : VITALDELAYTYPE01Z 	 := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
	tpd_A0_S0		 : VITALDELAYTYPE01 	 := (1.8 ns, 1.8 ns);
	tpd_B0_S0		 : VITALDELAYTYPE01 	 := (1.8 ns, 1.8 ns);
	tpd_CIN_S0		 : VITALDELAYTYPE01 	 := (1.8 ns, 1.8 ns);
	tpd_AS_S0		 : VITALDELAYTYPE01 	 := (1.8 ns, 1.8 ns);
	tpd_A0_COUT		 : VITALDELAYTYPE01 	 := (1.8 ns, 1.8 ns);
	tpd_B0_COUT		 : VITALDELAYTYPE01 	 := (1.8 ns, 1.8 ns);
	tpd_AS_COUT		 : VITALDELAYTYPE01 	 := (1.8 ns, 1.8 ns);
	tpd_CIN_COUT		 : VITALDELAYTYPE01 	 := (1.8 ns, 1.8 ns)
	);

PORT    (
	S0			 : OUT   std_logic;
	COUT			 : OUT   std_logic;
	A0			 : IN    std_logic := 'U';
	B0			 : IN    std_logic := 'U';
	CIN			 : IN    std_logic := 'U';
	AS			 : IN    std_logic := 'U'
	);

ATTRIBUTE VITAL_LEVEL0 OF CCU_AS : ENTITY IS TRUE ;

END CCU_AS;

-----------------------------------------------------------------------------
-- ARCHITECTURE declaration
-----------------------------------------------------------------------------
ARCHITECTURE VITAL_VF OF CCU_AS  IS
	ATTRIBUTE VITAL_LEVEL1 OF VITAL_VF : ARCHITECTURE IS TRUE;

	SIGNAL	A0_ipd			 : std_logic         := 'X';
	SIGNAL	B0_ipd			 : std_logic         := 'X';
	SIGNAL	CIN_ipd			 : std_logic         := 'X';
	SIGNAL	AS_ipd			 : std_logic         := 'X';
BEGIN
-----------------------------------------------------------------------------
-- INPUT PATH DELAYs
-----------------------------------------------------------------------------
WIREDELAY : BLOCK
BEGIN
	VitalWireDelay( A0_ipd, A0, tipd_A0 );
	VitalWireDelay( B0_ipd, B0, tipd_B0 );
	VitalWireDelay( CIN_ipd, CIN, tipd_CIN );
	VitalWireDelay( AS_ipd, AS, tipd_AS );
END BLOCK;

-----------------------------------------------------------------------------
-- Behavior Section
-----------------------------------------------------------------------------

VitalBehaviour_0 : PROCESS(A0_ipd,CIN_ipd,AS_ipd,B0_ipd)

VARIABLE 	S0_zd			 : std_ulogic;
VARIABLE 	out_1_zd		 : std_ulogic;
VARIABLE 	out_2_zd		 : std_ulogic;
VARIABLE 	out_3_zd		 : std_ulogic;
VARIABLE 	out_4_zd		 : std_ulogic;
VARIABLE 	COUT_zd			 : std_ulogic;
VARIABLE 	S0GLITCH_DATA		 : VitalGlitchDataType;
VARIABLE 	COUTGLITCH_DATA		 : VitalGlitchDataType;


BEGIN


--Functionality Section

out_1_zd	 := VitalXNOR2(AS_ipd,B0_ipd);
out_2_zd	 := VitalOR2(CIN_ipd,A0_ipd);
out_3_zd	 := VitalAND2(out_1_zd,out_2_zd);
out_4_zd	 := VitalAND2(CIN_ipd,A0_ipd);
COUT_zd		 := VitalOR2(out_4_zd,out_3_zd);
S0_zd		 := VitalXOR3(A0_ipd,CIN_ipd,out_1_zd);

--PathDelay Section

 VitalPathDelay01 ( S0, S0GLITCH_DATA, "S0", S0_zd,
	Paths => (
	0 => ( A0_ipd'LAST_EVENT, tpd_A0_S0, TRUE ),
	1 => ( B0_ipd'LAST_EVENT, tpd_B0_S0, TRUE ),
	2 => ( CIN_ipd'LAST_EVENT, tpd_CIN_S0, TRUE ),
	3 => ( AS_ipd'LAST_EVENT, tpd_AS_S0, TRUE ) ),
	DefaultDelay=>VitalZeroDelay01,
	Mode=>VitalInertial,
	XON=>TRUE,
	MsgOn=>TRUE,
	MsgSeverity=>WARNING );

 VitalPathDelay01 ( COUT, COUTGLITCH_DATA, "COUT", COUT_zd,
	Paths => (
	0 => ( A0_ipd'LAST_EVENT, tpd_A0_COUT, TRUE ),
	1 => ( B0_ipd'LAST_EVENT, tpd_B0_COUT, TRUE ),
	2 => ( AS_ipd'LAST_EVENT, tpd_AS_COUT, TRUE ),
	3 => ( CIN_ipd'LAST_EVENT, tpd_CIN_COUT, TRUE ) ),
	DefaultDelay=>VitalZeroDelay01,
	Mode=>VitalInertial,
	XON=>TRUE,
	MsgOn=>TRUE,
	MsgSeverity=>WARNING );


END PROCESS VitalBehaviour_0;


END VITAL_VF;
configuration CFG_CCU_AS_VITAL of CCU_AS is 
        for VITAL_VF
        end for; 
end CFG_CCU_AS_VITAL;
---------------------------------------------------------------------------------
-- VITAL model for cell CCU_DCP
---------------------------------------------------------------------------------
LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.VITAL_timing.all;
USE IEEE.VITAL_primitives.all;
LIBRARY VF1;
USE VF1.all;
USE VF1.VLOGTOVITAL_TABLES.all;
-----------------------------------------------------------------------------
--ENTITY DECLARATION
-----------------------------------------------------------------------------
ENTITY CCU_DCP IS

GENERIC (
	tipd_D			 : VITALDELAYTYPE01Z 	 := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
	tipd_LOAD		 : VITALDELAYTYPE01Z 	 := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
	tipd_CLK		 : VITALDELAYTYPE01Z 	 := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
	tipd_R			 : VITALDELAYTYPE01Z 	 := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
	tipd_S			 : VITALDELAYTYPE01Z 	 := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
	tipd_CIN		 : VITALDELAYTYPE01Z 	 := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
	tpd_CIN_COUT		 : VITALDELAYTYPE01 	 := (1 ns, 1 ns);
	tpd_R_Q			 : VITALDELAYTYPE01 	 := (1.44 ns, 1.44 ns);
	tpd_S_Q			 : VITALDELAYTYPE01 	 := (1.44 ns, 1.44 ns);
	tpd_CLK_Q		 : VITALDELAYTYPE01 	 := (1.44 ns, 1.44 ns);
	tpd_LOAD_Q		 : VITALDELAYTYPE01 	 := (2.69 ns, 2.69 ns);
	tpd_LOAD_COUT		 : VITALDELAYTYPE01 	 := (3.69 ns, 3.69 ns);
	tpd_D_Q			 : VITALDELAYTYPE01 	 := (2.69 ns, 2.69 ns);
	tpd_D_COUT		 : VITALDELAYTYPE01 	 := (3.69 ns, 3.69 ns)
	);

PORT    (
	Q			 : OUT   std_logic;
	COUT			 : OUT   std_logic;
	D			 : IN    std_logic := 'U';
	LOAD			 : IN    std_logic := 'U';
	CLK			 : IN    std_logic := 'U';
	R			 : IN    std_logic := 'U';
	S			 : IN    std_logic := 'U';
	CIN			 : IN    std_logic := 'U'
	);

ATTRIBUTE VITAL_LEVEL0 OF CCU_DCP : ENTITY IS TRUE ;

END CCU_DCP;

-----------------------------------------------------------------------------
-- ARCHITECTURE declaration
-----------------------------------------------------------------------------
ARCHITECTURE VITAL_VF OF CCU_DCP  IS
	ATTRIBUTE VITAL_LEVEL1 OF VITAL_VF : ARCHITECTURE IS TRUE;

	SIGNAL	Q_sig			 : std_logic         := 'X';
	SIGNAL	D_ipd			 : std_logic         := 'X';
	SIGNAL	LOAD_ipd		 : std_logic         := 'X';
	SIGNAL	CLK_ipd			 : std_logic         := 'X';
	SIGNAL	R_ipd			 : std_logic         := 'X';
	SIGNAL	S_ipd			 : std_logic         := 'X';
	SIGNAL	CIN_ipd			 : std_logic         := 'X';
	SIGNAL	Q_reg			 : std_logic         := 'X';
BEGIN
-----------------------------------------------------------------------------
-- INPUT PATH DELAYs
-----------------------------------------------------------------------------
WIREDELAY : BLOCK
BEGIN
	VitalWireDelay( D_ipd, D, tipd_D );
	VitalWireDelay( LOAD_ipd, LOAD, tipd_LOAD );
	VitalWireDelay( CLK_ipd, CLK, tipd_CLK );
	VitalWireDelay( R_ipd, R, tipd_R );
	VitalWireDelay( S_ipd, S, tipd_S );
	VitalWireDelay( CIN_ipd, CIN, tipd_CIN );
END BLOCK;

-----------------------------------------------------------------------------
-- Behavior Section
-----------------------------------------------------------------------------
VitalBehaviour_0 : PROCESS(LOAD_ipd,D_ipd,CLK_ipd,R_ipd,S_ipd,CIN_ipd,Q_sig)

VARIABLE 	load_zd			 : std_ulogic;
VARIABLE 	R_inv			 : std_ulogic;
VARIABLE 	S_inv			 : std_ulogic;
VARIABLE 	din0_zd			 : std_ulogic;
VARIABLE 	din1_zd			 : std_ulogic;
VARIABLE 	I1_zd			 : std_ulogic;
VARIABLE 	DIN_zd			 : std_ulogic;
VARIABLE 	Q_int_zd		 : std_ulogic;
VARIABLE 	notifier_zd		 : std_ulogic;
VARIABLE 	PrevDataIn0		 : std_logic_vector (0 to 3) ;
VARIABLE 	Q_zd			 : std_ulogic;
VARIABLE 	Q_reg_zd		 : std_ulogic;
VARIABLE 	O_zd			 : std_ulogic;
VARIABLE 	O1_zd			 : std_ulogic;
VARIABLE 	COUT_zd			 : std_ulogic;
VARIABLE 	Q_reg_tri		 : std_ulogic;
VARIABLE 	Bool_Condition01	 : BOOLEAN;
VARIABLE 	QGLITCH_DATA		 : VitalGlitchDataType;
VARIABLE 	COUTGLITCH_DATA		 : VitalGlitchDataType;
VARIABLE 	QsigGLITCH_DATA		 : VitalGlitchDataType;


BEGIN


--Functionality Section

load_zd		 := VitalINV(LOAD_ipd);
R_inv		 := VitalINV(R_ipd);
S_inv		 := VitalINV(S_ipd);
din0_zd		 := VitalAND2(LOAD_ipd,D_ipd);
notifier_zd	 := 'X';
I1_zd		 := VitalXNOR2(CIN_ipd,Q_sig);
O_zd		 := VitalOR2(Q_sig,CIN_ipd);
O1_zd		 := VitalAND2(load_zd,O_zd);
COUT_zd		 := VitalOR2(LOAD_ipd,O1_zd);
Q_reg_tri	 := Q_reg_zd;
din1_zd		 := VitalAND2(load_zd,I1_zd);
DIN_zd		 := VitalOR2(din0_zd,din1_zd);
VitalStateTable(
StateTable => dfftab,
DataIn => std_logic_vector'((DIN_zd),(CLK_ipd),(R_inv),(S_inv)),
Result => Q_int_zd,
PreviousDataIn => PrevDataIn0);
Q_reg_zd         :=Q_int_zd;
--Bool_Condition01 := (Q_int_zd /= ( not( '1')));
--Q_reg_zd	 := REG(Bool_Condition01,Q_int_zd);
--Q_reg_zd	 := TRIREG(Q_reg_zd,Q_reg_tri);
Q_zd		 := VitalBUF(Q_reg_zd);

--PathDelay Section

 VitalPathDelay01 ( Q, QGLITCH_DATA, "Q", Q_zd,
	Paths => (
	0 => ( R_ipd'LAST_EVENT, tpd_R_Q, TRUE ),
	1 => ( S_ipd'LAST_EVENT, tpd_S_Q, TRUE ),
	2 => ( CLK_ipd'LAST_EVENT, tpd_CLK_Q, TRUE ),
	3 => ( LOAD_ipd'LAST_EVENT, tpd_LOAD_Q, TRUE ),
	4 => ( D_ipd'LAST_EVENT, tpd_D_Q, TRUE ) ),
	DefaultDelay=>VitalZeroDelay01,
	Mode=>VitalInertial,
	XON=>TRUE,
	MsgOn=>TRUE,
	MsgSeverity=>WARNING );

 VitalPathDelay01 ( COUT, COUTGLITCH_DATA, "COUT", COUT_zd,
	Paths => (
	0 => ( CIN_ipd'LAST_EVENT, tpd_CIN_COUT, TRUE ),
	1 => ( LOAD_ipd'LAST_EVENT, tpd_LOAD_COUT, TRUE ),
	2 => ( D_ipd'LAST_EVENT, tpd_D_COUT, TRUE ) ),
	DefaultDelay=>VitalZeroDelay01,
	Mode=>VitalInertial,
	XON=>TRUE,
	MsgOn=>TRUE,
	MsgSeverity=>WARNING );

 VitalPathDelay01 ( Q_sig, QsigGLITCH_DATA, "Q_sig", Q_zd,
        Paths => (
        0 => ( 0.0 ns, (0.0 ns, 0.0 ns), FALSE  ) ),
        DefaultDelay=>VitalZeroDelay01,
        Mode=>VitalInertial,
        XON=>TRUE,
        MsgOn=>TRUE,
        MsgSeverity=>WARNING );
 
 


END PROCESS VitalBehaviour_0;


END VITAL_VF;
configuration CFG_CCU_DCP_VITAL of CCU_DCP is 
        for VITAL_VF
        end for; 
end CFG_CCU_DCP_VITAL;
---------------------------------------------------------------------------------
-- VITAL model for cell CCU_UCP
---------------------------------------------------------------------------------
LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.VITAL_timing.all;
USE IEEE.VITAL_primitives.all;
LIBRARY VF1;
USE VF1.all;
USE VF1.VLOGTOVITAL_TABLES.all;
-----------------------------------------------------------------------------
--ENTITY DECLARATION
-----------------------------------------------------------------------------
ENTITY CCU_UCP IS

GENERIC (
	tipd_D			 : VITALDELAYTYPE01Z 	 := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
	tipd_LOAD		 : VITALDELAYTYPE01Z 	 := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
	tipd_CLK		 : VITALDELAYTYPE01Z 	 := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
	tipd_R			 : VITALDELAYTYPE01Z 	 := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
	tipd_S			 : VITALDELAYTYPE01Z 	 := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
	tipd_CIN		 : VITALDELAYTYPE01Z 	 := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
	tpd_CIN_COUT		 : VITALDELAYTYPE01 	 := (1 ns, 1 ns);
	tpd_R_Q			 : VITALDELAYTYPE01 	 := (1.44 ns, 1.44 ns);
	tpd_S_Q			 : VITALDELAYTYPE01 	 := (1.44 ns, 1.44 ns);
	tpd_CLK_Q		 : VITALDELAYTYPE01 	 := (1.44 ns, 1.44 ns);
	tpd_LOAD_Q		 : VITALDELAYTYPE01 	 := (2.69 ns, 2.69 ns);
	tpd_LOAD_COUT		 : VITALDELAYTYPE01 	 := (3.69 ns, 3.69 ns);
	tpd_D_Q			 : VITALDELAYTYPE01 	 := (2.69 ns, 2.69 ns);
	tpd_D_COUT		 : VITALDELAYTYPE01 	 := (3.69 ns, 3.69 ns)
	);

PORT    (
	Q			 : OUT   std_logic;
	COUT			 : OUT   std_logic;
	D			 : IN    std_logic := 'U';
	LOAD			 : IN    std_logic := 'U';
	CLK			 : IN    std_logic := 'U';
	R			 : IN    std_logic := 'U';
	S			 : IN    std_logic := 'U';
	CIN			 : IN    std_logic := 'U'
	);

ATTRIBUTE VITAL_LEVEL0 OF CCU_UCP : ENTITY IS TRUE ;

END CCU_UCP;

-----------------------------------------------------------------------------
-- ARCHITECTURE declaration
-----------------------------------------------------------------------------
ARCHITECTURE VITAL_VF OF CCU_UCP  IS
	ATTRIBUTE VITAL_LEVEL1 OF VITAL_VF : ARCHITECTURE IS TRUE;

	SIGNAL	D_ipd			 : std_logic         := 'X';
	SIGNAL	LOAD_ipd		 : std_logic         := 'X';
	SIGNAL	CLK_ipd			 : std_logic         := 'X';
	SIGNAL	R_ipd			 : std_logic         := 'X';
	SIGNAL	S_ipd			 : std_logic         := 'X';
	SIGNAL	CIN_ipd			 : std_logic         := 'X';
	SIGNAL	Q_sig			 : std_logic         := 'X';
BEGIN
-----------------------------------------------------------------------------
-- INPUT PATH DELAYs
-----------------------------------------------------------------------------
WIREDELAY : BLOCK
BEGIN
	VitalWireDelay( D_ipd, D, tipd_D );
	VitalWireDelay( LOAD_ipd, LOAD, tipd_LOAD );
	VitalWireDelay( CLK_ipd, CLK, tipd_CLK );
	VitalWireDelay( R_ipd, R, tipd_R );
	VitalWireDelay( S_ipd, S, tipd_S );
	VitalWireDelay( CIN_ipd, CIN, tipd_CIN );
END BLOCK;

-----------------------------------------------------------------------------
-- Behavior Section
-----------------------------------------------------------------------------

VitalBehaviour_0 : PROCESS(Q_sig,LOAD_ipd,D_ipd,CLK_ipd,R_ipd,S_ipd,CIN_ipd)

VARIABLE 	load_zd			 : std_ulogic;
VARIABLE 	R_inverted			 : std_ulogic;
VARIABLE 	S_inverted			 : std_ulogic;
VARIABLE 	din0_zd			 : std_ulogic;
VARIABLE 	din1_zd			 : std_ulogic;
VARIABLE 	I1_zd			 : std_ulogic;
VARIABLE 	DIN_zd			 : std_ulogic;
VARIABLE 	Q_int_zd		 : std_ulogic;
VARIABLE 	notifier_zd		 : std_ulogic;
VARIABLE 	PrevDataIn0		 : std_logic_vector (0 to 3) ;
VARIABLE 	Q_zd			 : std_ulogic;
VARIABLE 	Q_reg_zd		 : std_ulogic;
VARIABLE 	COUT_zd			 : std_ulogic;
VARIABLE 	QGLITCH_DATA		 : VitalGlitchDataType;
VARIABLE 	QsigGLITCH_DATA		 : VitalGlitchDataType;
VARIABLE 	COUTGLITCH_DATA		 : VitalGlitchDataType;


BEGIN


--Functionality Section

load_zd		 := VitalINV(LOAD_ipd);
R_inverted		 := VitalINV(R_ipd);
S_inverted		 := VitalINV(S_ipd);
din0_zd		 := VitalAND2(LOAD_ipd,D_ipd);
notifier_zd	 := 'X';
Q_zd		 := VitalBUF(Q_sig);
I1_zd		 := VitalXOR2(CIN_ipd,Q_sig);
COUT_zd		 := VitalAND3(CIN_ipd,Q_sig,load_zd);
din1_zd		 := VitalAND2(load_zd,I1_zd);
DIN_zd		 := VitalOR2(din0_zd,din1_zd);
VitalStateTable(
StateTable => dfftab,
DataIn => std_logic_vector'((DIN_zd),(CLK_ipd),(R_inverted),(S_inverted)),
Result => Q_int_zd	,
PreviousDataIn => PrevDataIn0);

Q_reg_zd	 := Q_int_zd;


--PathDelay Section

 VitalPathDelay01 ( Q, QGLITCH_DATA, "Q", Q_zd,
	Paths => (
	0 => ( R_ipd'LAST_EVENT, tpd_R_Q, TRUE ),
	1 => ( S_ipd'LAST_EVENT, tpd_S_Q, TRUE ),
	2 => ( CLK_ipd'LAST_EVENT, tpd_CLK_Q, TRUE ),
	3 => ( LOAD_ipd'LAST_EVENT, tpd_LOAD_Q, TRUE ),
	4 => ( D_ipd'LAST_EVENT, tpd_D_Q, TRUE ) ),
	DefaultDelay=>VitalZeroDelay01,
	Mode=>VitalInertial,
	XON=>TRUE,
	MsgOn=>TRUE,
	MsgSeverity=>WARNING );

 VitalPathDelay01 ( COUT, COUTGLITCH_DATA, "COUT", COUT_zd,
	Paths => (
	0 => ( CIN_ipd'LAST_EVENT, tpd_CIN_COUT, TRUE ),
	1 => ( LOAD_ipd'LAST_EVENT, tpd_LOAD_COUT, TRUE ),
	2 => ( D_ipd'LAST_EVENT, tpd_D_COUT, TRUE ) ),
	DefaultDelay=>VitalZeroDelay01,
	Mode=>VitalInertial,
	XON=>TRUE,
	MsgOn=>TRUE,
	MsgSeverity=>WARNING );

 VitalPathDelay01 ( Q_sig, QsigGLITCH_DATA, "Q_sig", Q_reg_zd,
        Paths => (
        0 => ( 0.0 ns, (0.0 ns, 0.0 ns), FALSE  ) ),
        DefaultDelay=>VitalZeroDelay01,
        Mode=>VitalInertial,
        XON=>TRUE,
        MsgOn=>TRUE,
        MsgSeverity=>WARNING );
 



END PROCESS VitalBehaviour_0;


END VITAL_VF;
configuration CFG_CCU_UCP_VITAL of CCU_UCP is 
        for VITAL_VF
        end for; 
end CFG_CCU_UCP_VITAL;
---------------------------------------------------------------------------------
-- VITAL model for cell CCU_UDC
---------------------------------------------------------------------------------
LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.VITAL_timing.all;
USE IEEE.VITAL_primitives.all;
LIBRARY VF1;
USE VF1.all;
USE VF1.VLOGTOVITAL_TABLES.all;
-----------------------------------------------------------------------------
--ENTITY DECLARATION
-----------------------------------------------------------------------------
ENTITY CCU_UDC IS

GENERIC (
	tipd_UD			 : VITALDELAYTYPE01Z 	 := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
	tipd_CLK		 : VITALDELAYTYPE01Z 	 := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
	tipd_R			 : VITALDELAYTYPE01Z 	 := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
	tipd_S			 : VITALDELAYTYPE01Z 	 := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
	tipd_CIN		 : VITALDELAYTYPE01Z 	 := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
	TimingChecksOn           : BOOLEAN               := TRUE;
	ticd_CLK		 : VITALDELAYTYPE 	 := 0 ns;
	Xon                      : BOOLEAN               := FALSE;
	InstancePath             : STRING                := "*";
	MsgOn                    : BOOLEAN               := TRUE;
	tpw_CLK_posedge : VITALDELAYTYPE 	 := 4.4 ns;
	tpw_CLK_negedge : VITALDELAYTYPE 	 := 0 ns;
	tperiod_CLK_posedge : VITALDELAYTYPE 	 := 8.8 ns;
	ticd_R			 : VITALDELAYTYPE 	 := 0 ns;
	trecovery_CLK_R_posedge_posedge : VITALDELAYTYPE 	 := 2.2 ns;
	tremoval_CLK_R_posedge_posedge : VITALDELAYTYPE 	 := 0 ns;
	thold_R_CLK_posedge_posedge : VITALDELAYTYPE 	 := 2.2 ns;
	thold_R_CLK_negedge_posedge : VITALDELAYTYPE 	 := 0 ns;
	tsetup_R_CLK_noedge_posedge : VITALDELAYTYPE 	 := 0 ns;
	ticd_S			 : VITALDELAYTYPE 	 := 0 ns;
	trecovery_CLK_S_posedge_posedge : VITALDELAYTYPE 	 := 2.2 ns;
	tremoval_CLK_S_posedge_posedge : VITALDELAYTYPE 	 := 0 ns;
	thold_S_CLK_posedge_posedge : VITALDELAYTYPE 	 := 2.2 ns;
	thold_S_CLK_negedge_posedge : VITALDELAYTYPE 	 := 0 ns;
	tsetup_S_CLK_noedge_posedge : VITALDELAYTYPE 	 := 0 ns;
	tpd_CIN_COUT		 : VITALDELAYTYPE01 	 := (1 ns, 1 ns);
	tpd_UD_COUT		 : VITALDELAYTYPE01 	 := (1 ns, 1 ns);
	tpd_UD_Q		 : VITALDELAYTYPE01 	 := (2.44 ns, 2.44 ns);
	tpd_CIN_Q		 : VITALDELAYTYPE01 	 := (2.44 ns, 2.44 ns);
	tpd_CLK_Q		 : VITALDELAYTYPE01 	 := (1.44 ns, 1.44 ns);
	tpd_R_Q			 : VITALDELAYTYPE01 	 := (1.44 ns, 1.44 ns);
	tpd_S_Q			 : VITALDELAYTYPE01 	 := (1.44 ns, 1.44 ns)
	);

PORT    (
	Q			 : OUT   std_logic;
	COUT			 : OUT   std_logic;
	UD			 : IN    std_logic := 'U';
	CLK			 : IN    std_logic := 'U';
	R			 : IN    std_logic := 'U';
	S			 : IN    std_logic := 'U';
	CIN			 : IN    std_logic := 'U'
	);

ATTRIBUTE VITAL_LEVEL0 OF CCU_UDC : ENTITY IS TRUE ;

END CCU_UDC;

-----------------------------------------------------------------------------
-- ARCHITECTURE declaration
-----------------------------------------------------------------------------
ARCHITECTURE VITAL_VF OF CCU_UDC  IS
	ATTRIBUTE VITAL_LEVEL1 OF VITAL_VF : ARCHITECTURE IS TRUE;

	SIGNAL	UD_ipd			 : std_logic         := 'X';
	SIGNAL	CLK_ipd			 : std_logic         := 'X';
	SIGNAL	R_ipd			 : std_logic         := 'X';
	SIGNAL	S_ipd			 : std_logic         := 'X';
	SIGNAL	CIN_ipd			 : std_logic         := 'X';
	SIGNAL	CLK_dly			 : std_ulogic        := 'X';
	SIGNAL	R_dly			 : std_ulogic        := 'X';
	SIGNAL	S_dly			 : std_ulogic        := 'X';
	SIGNAL	Q_sig			 : std_ulogic        := 'X';
BEGIN
-----------------------------------------------------------------------------
-- INPUT PATH DELAYs
-----------------------------------------------------------------------------
WIREDELAY : BLOCK
BEGIN
	VitalWireDelay( UD_ipd, UD, tipd_UD );
	VitalWireDelay( CLK_ipd, CLK, tipd_CLK );
	VitalWireDelay( R_ipd, R, tipd_R );
	VitalWireDelay( S_ipd, S, tipd_S );
	VitalWireDelay( CIN_ipd, CIN, tipd_CIN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
	VitalSignalDelay ( CLK_dly, CLK_ipd, ticd_CLK);
	VitalSignalDelay ( R_dly, R_ipd, ticd_R);
	VitalSignalDelay ( S_dly, S_ipd, ticd_S);
END BLOCK;

-----------------------------------------------------------------------------
-- Behavior Section
-----------------------------------------------------------------------------

VitalBehaviour_0 : PROCESS(Q_sig,R_ipd,S_ipd,R_dly,UD_ipd,CIN_ipd,CLK_dly,S_dly)

VARIABLE 	Tviol_CLK_flag1		 : std_ulogic		 := '0';
VARIABLE 	PeriodData_CLK1		 : VitalPeriodDataType	 := VitalPeriodDataInit;
VARIABLE 	Tviol_CLK_flag2		 : std_ulogic		 := '0';
VARIABLE 	PeriodData_CLK2		 : VitalPeriodDataType	 := VitalPeriodDataInit;
VARIABLE 	Tviol_R_CLK_flag3	 : std_ulogic		 := '0';
VARIABLE 	TimingData_CLK_R3	 : VitalTimingDataType	 := VitalTimingDataInit;
VARIABLE 	Tviol_CLK_R_flag4	 : std_ulogic		 := '0';
VARIABLE 	TimingData_R_CLK4	 : VitalTimingDataType	 := VitalTimingDataInit;
VARIABLE 	Tviol_S_CLK_flag5	 : std_ulogic		 := '0';
VARIABLE 	TimingData_CLK_S5	 : VitalTimingDataType	 := VitalTimingDataInit;
VARIABLE 	Tviol_CLK_S_flag6	 : std_ulogic		 := '0';
VARIABLE 	TimingData_S_CLK6	 : VitalTimingDataType	 := VitalTimingDataInit;
VARIABLE 	ud_zd			 : std_ulogic;
VARIABLE 	S0_zd			 : std_ulogic;
VARIABLE 	A0_zd			 : std_ulogic;
VARIABLE 	c0_zd			 : std_ulogic;
VARIABLE 	c1_zd			 : std_ulogic;
VARIABLE 	c2_zd			 : std_ulogic;
VARIABLE 	COUT_zd			 : std_ulogic;
VARIABLE 	Q_int_zd		 : std_ulogic;
VARIABLE 	R_inverted		 : std_ulogic;
VARIABLE 	S_inverted		 : std_ulogic;
VARIABLE 	notifier_zd		 : std_ulogic;
VARIABLE 	PrevDataIn0		 : std_logic_vector (0 to 3) ;
VARIABLE 	Q_reg_zd		 : std_ulogic;
VARIABLE 	Q_zd			 : std_ulogic;
VARIABLE 	R_S_zd			 : std_ulogic;
VARIABLE 	QGLITCH_DATA		 : VitalGlitchDataType;
VARIABLE 	COUTGLITCH_DATA		 : VitalGlitchDataType;
VARIABLE 	QsigGLITCH_DATA		 : VitalGlitchDataType;
VARIABLE 	Violation_Flag		 : std_ulogic;


BEGIN

--Timing Check Section

IF(TimingChecksOn) THEN
VitalPeriodPulseCheck(Violation => Tviol_CLK_flag1,
PeriodData => PeriodData_CLK1,
TestSignal => CLK_dly,
TestSignalName => "CLK",
TestDelay => 0 ns,
Period => 0 ns,
PulseWidthHigh => tpw_CLK_posedge,
PulseWidthLow => tpw_CLK_negedge,
CheckEnabled => ( To_X01( R_S_zd )= '1' ),
HeaderMsg => InstancePath & "/CCU_UDC",
Xon => Xon,
MsgOn => MsgOn,
MsgSeverity => WARNING);


VitalPeriodPulseCheck(Violation => Tviol_CLK_flag2,
PeriodData => PeriodData_CLK2,
TestSignal => CLK_dly,
TestSignalName => "CLK",
TestDelay => 0 ns,
Period => tperiod_CLK_posedge,
PulseWidthHigh => 0 ns,
PulseWidthLow => 0 ns,
CheckEnabled => posedge( CLK_dly'LAST_VALUE, CLK_dly ) AND ( To_X01( R_S_zd )= '1' ),
HeaderMsg => InstancePath & "/CCU_UDC",
Xon => Xon,
MsgOn => MsgOn,
MsgSeverity => WARNING);


VitalRecoveryRemovalCheck(Violation => Tviol_R_CLK_flag3,
TimingData => TimingData_CLK_R3,
TestSignal => CLK_dly,
TestSignalName => "CLK",
TestDelay => 0 ns,
RefSignal => R_dly,
RefSignalName => "R",
RefDelay => 0 ns,
Recovery => trecovery_CLK_R_posedge_posedge,
Removal => tremoval_CLK_R_posedge_posedge,
ActiveLow => FALSE,
CheckEnabled => ( To_X01( S_ipd )= '0' ),
RefTransition => '/',
HeaderMsg =>InstancePath & "/CCU_UDC",
Xon => Xon,
MsgOn => MsgOn,
MsgSeverity => WARNING);


VitalSetupHoldCheck(Violation => Tviol_CLK_R_flag4,
TimingData => TimingData_R_CLK4,
TestSignal => R_dly,
TestSignalName => "R",
TestDelay => 0 ns,
RefSignal => CLK_dly,
RefSignalName => "CLK",
RefDelay => 0 ns,
SetupHigh => tsetup_R_CLK_noedge_posedge,
SetupLow => tsetup_R_CLK_noedge_posedge,
HoldHigh => thold_R_CLK_posedge_posedge,
HoldLow => thold_R_CLK_negedge_posedge,
CheckEnabled => ( To_X01( S_ipd )= '0' ),
RefTransition => '/',
HeaderMsg => InstancePath & "/CCU_UDC",
Xon => Xon,
MsgOn => MsgOn,
MsgSeverity => WARNING);


VitalRecoveryRemovalCheck(Violation => Tviol_S_CLK_flag5,
TimingData => TimingData_CLK_S5,
TestSignal => CLK_dly,
TestSignalName => "CLK",
TestDelay => 0 ns,
RefSignal => S_dly,
RefSignalName => "S",
RefDelay => 0 ns,
Recovery => trecovery_CLK_S_posedge_posedge,
Removal => tremoval_CLK_S_posedge_posedge,
ActiveLow => FALSE,
CheckEnabled => ( To_X01( R_dly )= '0' ),
RefTransition => '/',
HeaderMsg =>InstancePath & "/CCU_UDC",
Xon => Xon,
MsgOn => MsgOn,
MsgSeverity => WARNING);


VitalSetupHoldCheck(Violation => Tviol_CLK_S_flag6,
TimingData => TimingData_S_CLK6,
TestSignal => S_dly,
TestSignalName => "S",
TestDelay => 0 ns,
RefSignal => CLK_dly,
RefSignalName => "CLK",
RefDelay => 0 ns,
SetupHigh => tsetup_S_CLK_noedge_posedge,
SetupLow => tsetup_S_CLK_noedge_posedge,
HoldHigh => thold_S_CLK_posedge_posedge,
HoldLow => thold_S_CLK_negedge_posedge,
CheckEnabled => ( To_X01( R_dly )= '0' ),
RefTransition => '/',
HeaderMsg => InstancePath & "/CCU_UDC",
Xon => Xon,
MsgOn => MsgOn,
MsgSeverity => WARNING);


END IF;   -- Timing Check Section

--Functionality Section

Violation_Flag	 := (((((Tviol_CLK_flag1 or Tviol_CLK_flag2) or Tviol_R_CLK_flag3) or Tviol_CLK_R_flag4) or Tviol_S_CLK_flag5) or Tviol_CLK_S_flag6);
ud_zd		 := VitalINV(UD_ipd);
R_inverted		 := VitalINV(R_ipd);
S_inverted		 := VitalINV(S_ipd);
c2_zd		 := VitalAND2(ud_zd,CIN_ipd);
notifier_zd	 := 'X';
A0_zd		 := VitalBUF(Q_sig);
Q_zd		 := VitalBUF(Q_sig);
R_S_zd		 := VitalAND2(R_inverted,S_inverted);
S0_zd		 := VitalXOR3(A0_zd,ud_zd,CIN_ipd);
c0_zd		 := VitalAND2(A0_zd,ud_zd);
c1_zd		 := VitalAND2(A0_zd,CIN_ipd);
COUT_zd		 := VitalOR3(c0_zd,c1_zd,c2_zd);
VitalStateTable(
StateTable => dfftab,
DataIn => std_logic_vector'((S0_zd),(CLK_dly),(R_inverted),(S_inverted)),
Result => Q_int_zd	,
PreviousDataIn => PrevDataIn0);

Q_int_zd	 := (Violation_Flag xor Q_int_zd);
Q_reg_zd	 := Q_int_zd;

--PathDelay Section

 VitalPathDelay01 ( Q, QGLITCH_DATA, "Q", Q_zd,
	Paths => (
	0 => ( UD_ipd'LAST_EVENT, tpd_UD_Q, TRUE ),
	1 => ( CIN_ipd'LAST_EVENT, tpd_CIN_Q, TRUE ),
	2 => ( CLK_dly'LAST_EVENT, tpd_CLK_Q, TRUE ),
	3 => ( R_dly'LAST_EVENT, tpd_R_Q, TRUE ),
	4 => ( S_dly'LAST_EVENT, tpd_S_Q, TRUE ) ),
	DefaultDelay=>VitalZeroDelay01,
	Mode=>VitalInertial,
	XON=>TRUE,
	MsgOn=>TRUE,
	MsgSeverity=>WARNING );

 VitalPathDelay01 ( COUT, COUTGLITCH_DATA, "COUT", COUT_zd,
	Paths => (
	0 => ( CIN_ipd'LAST_EVENT, tpd_CIN_COUT, TRUE ),
	1 => ( UD_ipd'LAST_EVENT, tpd_UD_COUT, TRUE ) ),
	DefaultDelay=>VitalZeroDelay01,
	Mode=>VitalInertial,
	XON=>TRUE,
	MsgOn=>TRUE,
	MsgSeverity=>WARNING );

 VitalPathDelay01 ( Q_sig, QsigGLITCH_DATA, "Q_sig", Q_reg_zd,
        Paths => (
        0 => ( 0.0 ns, (0.0 ns, 0.0 ns), FALSE  ) ),
        DefaultDelay=>VitalZeroDelay01,
        Mode=>VitalInertial,
        XON=>TRUE,
        MsgOn=>TRUE,
        MsgSeverity=>WARNING );
 



END PROCESS VitalBehaviour_0;


END VITAL_VF;
configuration CFG_CCU_UDC_VITAL of CCU_UDC is 
        for VITAL_VF
        end for; 
end CFG_CCU_UDC_VITAL;
----- VITAL model for cell CLKI -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity CLKI is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_PAD_O                       :	VitalDelayType01 := (1.25 ns, 1.25 ns);
      tipd_PAD                        :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      PAD                             :	in    STD_ULOGIC;
      O                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of CLKI : entity is TRUE;
end CLKI;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library VF1;
architecture VITAL_VF of CLKI is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL PAD_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (PAD_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS O_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE O_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      O_zd := TO_X01(PAD_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => O,
       GlitchData => O_GlitchData,
       OutSignalName => "O",
       OutTemp => O_zd,
       Paths => (0 => (PAD_ipd'last_event, tpd_PAD_O, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;

configuration CFG_CLKI_VITAL of CLKI is 
        for VITAL_VF
        end for; 
end CFG_CLKI_VITAL;
----- VITAL model for cell COM_UDCP -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;
library VF1;
use VF1.all;


-- entity declaration --
entity COM_UDCP is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_LOAD_Q                     :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_CNTEN_Q                      :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_A_Q                        :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_UD_Q                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_CIN_Q                      :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_D_Q                        :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_LOAD_COUT                  :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_CNTEN_COUT                   :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_A_COUT                     :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_UD_COUT                    :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_CIN_COUT                   :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_LOAD                      :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CNTEN                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_UD                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CIN                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      LOAD                           :	in    STD_ULOGIC;
      CNTEN                            :	in    STD_ULOGIC;
      A                              :	in    STD_ULOGIC;
      UD                             :	in    STD_ULOGIC;
      CIN                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      COUT                           :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of COM_UDCP : entity is TRUE;
end COM_UDCP;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library VF1;
architecture VITAL_VF of COM_UDCP is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL LOAD_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CNTEN_ipd	 : STD_ULOGIC := 'X';
   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL UD_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CIN_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (LOAD_ipd, LOAD, tipd_LOAD);
   VitalWireDelay (CNTEN_ipd, CNTEN, tipd_CNTEN);
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (UD_ipd, UD, tipd_UD);
   VitalWireDelay (CIN_ipd, CIN, tipd_CIN);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, LOAD_ipd, CNTEN_ipd, A_ipd, UD_ipd, CIN_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);
   ALIAS COUT_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;
   VARIABLE COUT_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd :=
       ((((A_ipd) AND ((NOT CNTEN_ipd))) OR ((((NOT UD_ipd)) XOR (A_ipd) XOR
         (CIN_ipd)) AND (CNTEN_ipd))) AND ((NOT LOAD_ipd))) OR ((D_ipd) AND
         (LOAD_ipd));
      COUT_zd :=
       (CNTEN_ipd) AND ((NOT LOAD_ipd)) AND (((CIN_ipd) AND (A_ipd)) OR (((NOT
         UD_ipd)) AND (A_ipd)) OR (((NOT UD_ipd)) AND (CIN_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (LOAD_ipd'last_event, tpd_LOAD_Q, TRUE),
                 1 => (CNTEN_ipd'last_event, tpd_CNTEN_Q, TRUE),
                 2 => (A_ipd'last_event, tpd_A_Q, TRUE),
                 3 => (UD_ipd'last_event, tpd_UD_Q, TRUE),
                 4 => (CIN_ipd'last_event, tpd_CIN_Q, TRUE),
                 5 => (D_ipd'last_event, tpd_D_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);
      VitalPathDelay01 (
       OutSignal => COUT,
       GlitchData => COUT_GlitchData,
       OutSignalName => "COUT",
       OutTemp => COUT_zd,
       Paths => (0 => (LOAD_ipd'last_event, tpd_LOAD_COUT, TRUE),
                 1 => (CNTEN_ipd'last_event, tpd_CNTEN_COUT, TRUE),
                 2 => (A_ipd'last_event, tpd_A_COUT, TRUE),
                 3 => (UD_ipd'last_event, tpd_UD_COUT, TRUE),
                 4 => (CIN_ipd'last_event, tpd_CIN_COUT, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;

configuration CFG_COM_UDCP_VITAL of COM_UDCP is 
        for VITAL_VF
        end for; 
end CFG_COM_UDCP_VITAL;
----- VITAL model for cell DEMUX2 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DEMUX2 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_EN_O0                      :	VitalDelayType01 := (1.250 ns, 1.250 ns);
      tpd_S0_O0                      :	VitalDelayType01 := (1.250 ns, 1.250 ns);
      tpd_EN_O1                      :	VitalDelayType01 := (1.250 ns, 1.250 ns);
      tpd_S0_O1                      :	VitalDelayType01 := (1.250 ns, 1.250 ns);
      tipd_EN                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      EN                             :	in    STD_ULOGIC;
      S0                             :	in    STD_ULOGIC;
      O0                             :	out   STD_ULOGIC;
      O1                             :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DEMUX2 : entity is TRUE;
end DEMUX2;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library VF1;
architecture VITAL_VF of DEMUX2 is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL EN_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S0_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (EN_ipd, EN, tipd_EN);
   VitalWireDelay (S0_ipd, S0, tipd_S0);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (EN_ipd, S0_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS O0_zd : STD_LOGIC is Results(1);
   ALIAS O1_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE O0_GlitchData	: VitalGlitchDataType;
   VARIABLE O1_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      O0_zd := ((NOT S0_ipd)) AND (EN_ipd);
      O1_zd := (S0_ipd) AND (EN_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => O0,
       GlitchData => O0_GlitchData,
       OutSignalName => "O0",
       OutTemp => O0_zd,
       Paths => (0 => (EN_ipd'last_event, tpd_EN_O0, TRUE),
                 1 => (S0_ipd'last_event, tpd_S0_O0, TRUE)),
       Mode => VitalInertial,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);
      VitalPathDelay01 (
       OutSignal => O1,
       GlitchData => O1_GlitchData,
       OutSignalName => "O1",
       OutTemp => O1_zd,
       Paths => (0 => (EN_ipd'last_event, tpd_EN_O1, TRUE),
                 1 => (S0_ipd'last_event, tpd_S0_O1, TRUE)),
       Mode => VitalInertial,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;

configuration CFG_DEMUX2_VITAL of DEMUX2 is 
        for VITAL_VF
        end for; 
end CFG_DEMUX2_VITAL;
----- VITAL model for cell DEMUX4 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DEMUX4 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_EN_O0                      :	VitalDelayType01 := (1.25 ns, 1.25 ns);
      tpd_S0_O0                      :	VitalDelayType01 := (1.25 ns, 1.25 ns);
      tpd_S1_O0                      :	VitalDelayType01 := (1.25 ns, 1.25 ns);
      tpd_EN_O1                      :	VitalDelayType01 := (1.25 ns, 1.25 ns);
      tpd_S0_O1                      :	VitalDelayType01 := (1.25 ns, 1.25 ns);
      tpd_S1_O1                      :	VitalDelayType01 := (1.25 ns, 1.25 ns);
      tpd_EN_O2                      :	VitalDelayType01 := (1.25 ns, 1.25 ns);
      tpd_S0_O2                      :	VitalDelayType01 := (1.25 ns, 1.25 ns);
      tpd_S1_O2                      :	VitalDelayType01 := (1.25 ns, 1.25 ns);
      tpd_EN_O3                      :	VitalDelayType01 := (1.25 ns, 1.25 ns);
      tpd_S0_O3                      :	VitalDelayType01 := (1.25 ns, 1.25 ns);
      tpd_S1_O3                      :	VitalDelayType01 := (1.25 ns, 1.25 ns);
      tipd_EN                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      EN                             :	in    STD_ULOGIC;
      S0                             :	in    STD_ULOGIC;
      S1                             :	in    STD_ULOGIC;
      O0                             :	out   STD_ULOGIC;
      O1                             :	out   STD_ULOGIC;
      O2                             :	out   STD_ULOGIC;
      O3                             :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DEMUX4 : entity is TRUE;
end DEMUX4;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library VF1;
architecture VITAL_VF of DEMUX4 is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL EN_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S1_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (EN_ipd, EN, tipd_EN);
   VitalWireDelay (S0_ipd, S0, tipd_S0);
   VitalWireDelay (S1_ipd, S1, tipd_S1);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (EN_ipd, S0_ipd, S1_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 4) := (others => 'X');
   ALIAS O0_zd : STD_LOGIC is Results(1);
   ALIAS O1_zd : STD_LOGIC is Results(2);
   ALIAS O2_zd : STD_LOGIC is Results(3);
   ALIAS O3_zd : STD_LOGIC is Results(4);

   -- output glitch detection variables
   VARIABLE O0_GlitchData	: VitalGlitchDataType;
   VARIABLE O1_GlitchData	: VitalGlitchDataType;
   VARIABLE O2_GlitchData	: VitalGlitchDataType;
   VARIABLE O3_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      O0_zd := ((NOT S0_ipd)) AND (EN_ipd) AND ((NOT S1_ipd));
      O1_zd := (S0_ipd) AND (EN_ipd) AND ((NOT S1_ipd));
      O2_zd := ((NOT S0_ipd)) AND (EN_ipd) AND (S1_ipd);
      O3_zd := (S0_ipd) AND (EN_ipd) AND (S1_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => O0,
       GlitchData => O0_GlitchData,
       OutSignalName => "O0",
       OutTemp => O0_zd,
       Paths => (0 => (EN_ipd'last_event, tpd_EN_O0, TRUE),
                 1 => (S0_ipd'last_event, tpd_S0_O0, TRUE),
                 2 => (S1_ipd'last_event, tpd_S1_O0, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);
      VitalPathDelay01 (
       OutSignal => O1,
       GlitchData => O1_GlitchData,
       OutSignalName => "O1",
       OutTemp => O1_zd,
       Paths => (0 => (EN_ipd'last_event, tpd_EN_O1, TRUE),
                 1 => (S0_ipd'last_event, tpd_S0_O1, TRUE),
                 2 => (S1_ipd'last_event, tpd_S1_O1, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);
      VitalPathDelay01 (
       OutSignal => O2,
       GlitchData => O2_GlitchData,
       OutSignalName => "O2",
       OutTemp => O2_zd,
       Paths => (0 => (EN_ipd'last_event, tpd_EN_O2, TRUE),
                 1 => (S0_ipd'last_event, tpd_S0_O2, TRUE),
                 2 => (S1_ipd'last_event, tpd_S1_O2, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);
      VitalPathDelay01 (
       OutSignal => O3,
       GlitchData => O3_GlitchData,
       OutSignalName => "O3",
       OutTemp => O3_zd,
       Paths => (0 => (EN_ipd'last_event, tpd_EN_O3, TRUE),
                 1 => (S0_ipd'last_event, tpd_S0_O3, TRUE),
                 2 => (S1_ipd'last_event, tpd_S1_O3, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;

configuration CFG_DEMUX4_VITAL of DEMUX4 is 
        for VITAL_VF
        end for; 
end CFG_DEMUX4_VITAL;
----- VITAL model for cell DFF -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;

LIBRARY VF1 ;
use VF1.VLOGTOVITAL_TABLES.all;



-- entity declaration --
entity DFF is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_CLK_Q                      :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tsetup_D_CLK_noedge_posedge    :	VitalDelayType := 2.200 ns;
      thold_D_CLK_noedge_posedge     :	VitalDelayType := 2.200 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 8.800 ns;
      tpw_CLK_posedge                :	VitalDelayType := 4.400 ns;
      ticd_CLK                       :	VitalDelayType := 0.000 ns;
      tisd_D_CLK                     :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFF : entity is TRUE;
end DFF;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library VF1;
architecture VITAL_VF of DFF is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL D_CLK_dly	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   VitalSignalDelay (CLK_dly, CLK_ipd, ticd_CLK);
   VitalSignalDelay (D_CLK_dly, D_ipd, tisd_D_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (CLK_dly, D_CLK_dly)

   -- timing check results
   VARIABLE Tviol_D_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 3);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_posedge,
          TimingData              => Tmkr_D_CLK_posedge,
          TestSignal              => D_CLK_dly,
          TestSignalName          => "D",
          TestDelay               => tisd_D_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          SetupHigh               => tsetup_D_CLK_noedge_posedge,
          SetupLow                => tsetup_D_CLK_noedge_posedge,
          HoldHigh                => thold_D_CLK_noedge_posedge,
          HoldLow                 => thold_D_CLK_noedge_posedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFF",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_dly,
          TestSignalName          => "CLK",
          TestDelay               => ticd_CLK,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFF",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_posedge or Pviol_CLK;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => dfftab,
        DataIn => (
               D_CLK_dly, CLK_dly, '1','1'));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (CLK_dly'last_event, tpd_CLK_Q, TRUE)),
       Mode => VitalInertial,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;

configuration CFG_DFF_VITAL of DFF is 
        for VITAL_VF
        end for; 
end CFG_DFF_VITAL;
----- VITAL model for cell DFFC -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;

LIBRARY VF1 ;
use VF1.VLOGTOVITAL_TABLES.all;



-- entity declaration --
entity DFFC is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_CLK_Q                      :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tsetup_D_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      thold_D_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      tsetup_CE_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      thold_CE_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      tpw_CLK_posedge        :	VitalDelayType := 4.400 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 8.800 ns;
      ticd_CLK                       :	VitalDelayType := 0.000 ns;
      tisd_D_CLK                     :	VitalDelayType := 0.000 ns;
      tisd_CE_CLK                     :	VitalDelayType := 0.000 ns;
      tipd_CE                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      CE                             :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFFC : entity is TRUE;
end DFFC;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library VF1;
architecture VITAL_VF of DFFC is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL CE_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL D_CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL CE_CLK_dly	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (CE_ipd, CE, tipd_CE);
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   VitalSignalDelay (CLK_dly, CLK_ipd, ticd_CLK);
   VitalSignalDelay (D_CLK_dly, D_ipd, tisd_D_CLK);
   VitalSignalDelay (CE_CLK_dly, CE_ipd, tisd_CE_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (CE_ipd, CLK_dly, D_CLK_dly, CE_CLK_dly)

   -- timing check results
   VARIABLE Tviol_D_CLK_CE_EQ_1_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_CE_EQ_1_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CE_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CE_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK_CE_EQ_1	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK_CE_EQ_1	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 4);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_CE_EQ_1_posedge,
          TimingData              => Tmkr_D_CLK_CE_EQ_1_posedge,
          TestSignal              => D_CLK_dly,
          TestSignalName          => "D",
          TestDelay               => tisd_D_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          SetupHigh               => tsetup_D_CLK_noedge_posedge,
          SetupLow                => tsetup_D_CLK_noedge_posedge,
          HoldHigh                => thold_D_CLK_noedge_posedge,
          HoldLow                 => thold_D_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(CE_ipd) = '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFFC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);

         VitalSetupHoldCheck (
          Violation               => Tviol_CE_CLK_posedge,
          TimingData              => Tmkr_CE_CLK_posedge,
          TestSignal              => CE_CLK_dly,
          TestSignalName          => "CE",
          TestDelay               => tisd_CE_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          SetupHigh               => tsetup_CE_CLK_noedge_posedge,
          SetupLow                => tsetup_CE_CLK_noedge_posedge,
          HoldHigh                => thold_CE_CLK_noedge_posedge,
          HoldLow                 => thold_CE_CLK_noedge_posedge,
          CheckEnabled            => TRUE, 
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFFC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);

         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK_CE_EQ_1,
          PeriodData              => PInfo_CLK_CE_EQ_1,
          TestSignal              => CLK_dly,
          TestSignalName          => "CLK",
          TestDelay               => ticd_CLK,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
			TO_X01(CE_ipd) = '1',
          HeaderMsg               => InstancePath & "/DFFC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_CE_EQ_1_posedge or Tviol_CE_CLK_posedge or Pviol_CLK_CE_EQ_1;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => dffcetab,
        DataIn => (
               D_CLK_dly, CLK_dly,'1','1', CE_CLK_dly));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (CLK_dly'last_event, tpd_CLK_Q, TRUE)),
       Mode => VitalInertial,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;

configuration CFG_DFFC_VITAL of DFFC is 
        for VITAL_VF
        end for; 
end CFG_DFFC_VITAL;
----- VITAL model for cell DFFCR -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;

LIBRARY VF1 ;
use VF1.VLOGTOVITAL_TABLES.all;



-- entity declaration --
entity DFFCR is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_R_Q                        :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tsetup_D_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      thold_D_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      tsetup_CE_CLK_posedge_posedge :	VitalDelayType := 2.200 ns;
      thold_CE_CLK_posedge_posedge :	VitalDelayType := 2.200 ns;
      tpw_CLK_posedge :	VitalDelayType := 4.400 ns;
      tperiod_CLK_posedge :	VitalDelayType := 8.800 ns;
      trecovery_R_CLK_posedge_posedge :	VitalDelayType := 2.200 ns;
      thold_R_CLK_posedge_posedge :	VitalDelayType := 2.200 ns;
      ticd_CLK                       :	VitalDelayType := 0.000 ns;
      tisd_D_CLK                     :	VitalDelayType := 0.000 ns;
      tisd_CE_CLK                     :	VitalDelayType := 0.000 ns;
      tisd_R_CLK                     :	VitalDelayType := 0.000 ns;
      tipd_CE                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_R                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      CE                             :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      R                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFFCR : entity is TRUE;
end DFFCR;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library VF1;
architecture VITAL_VF of DFFCR is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL CE_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL R_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL D_CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL CE_CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL R_CLK_dly	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (CE_ipd, CE, tipd_CE);
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (R_ipd, R, tipd_R);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   VitalSignalDelay (CLK_dly, CLK_ipd, ticd_CLK);
   VitalSignalDelay (D_CLK_dly, D_ipd, tisd_D_CLK);
   VitalSignalDelay (CE_CLK_dly, CE_ipd, tisd_CE_CLK);
   VitalSignalDelay (R_CLK_dly, R_ipd, tisd_R_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (CE_ipd, CLK_dly, D_CLK_dly, R_CLK_dly, CE_CLK_dly)

   -- timing check results
   VARIABLE Tviol_D_CLK_CE_EQ_1_ANB_R_EQ_1_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_CE_EQ_1_ANB_R_EQ_1_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CE_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CE_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_R_CLK_CE_EQ_1_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_R_CLK_CE_EQ_1_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK_CE_EQ_1_ANB_R_EQ_1	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK_CE_EQ_1_ANB_R_EQ_1	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 4);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_CE_EQ_1_ANB_R_EQ_1_posedge,
          TimingData              => Tmkr_D_CLK_CE_EQ_1_ANB_R_EQ_1_posedge,
          TestSignal              => D_CLK_dly,
          TestSignalName          => "D",
          TestDelay               => tisd_D_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          SetupHigh               => tsetup_D_CLK_noedge_posedge,
          SetupLow                => tsetup_D_CLK_noedge_posedge,
          HoldHigh                => thold_D_CLK_noedge_posedge,
          HoldLow                 => thold_D_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((R_CLK_dly) AND (CE_ipd)) = '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFFCR",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_CE_CLK_posedge,
          TimingData              => Tmkr_CE_CLK_posedge,
          TestSignal              => CE_CLK_dly,
          TestSignalName          => "CE",
          TestDelay               => tisd_CE_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          SetupHigh               => tsetup_CE_CLK_posedge_posedge,
          SetupLow                => tsetup_CE_CLK_posedge_posedge,
          HoldHigh                => thold_CE_CLK_posedge_posedge,
          HoldLow                 => thold_CE_CLK_posedge_posedge,
          CheckEnabled            => TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFFCR",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_R_CLK_CE_EQ_1_posedge,
          TimingData              => Tmkr_R_CLK_CE_EQ_1_posedge,
          TestSignal              => R_CLK_dly,
          TestSignalName          => "R",
          TestDelay               => tisd_R_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          Recovery                => trecovery_R_CLK_posedge_posedge,
          Removal                 => thold_R_CLK_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TO_X01(CE_ipd) = '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFFCR",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK_CE_EQ_1_ANB_R_EQ_1,
          PeriodData              => PInfo_CLK_CE_EQ_1_ANB_R_EQ_1,
          TestSignal              => CLK_dly,
          TestSignalName          => "CLK",
          TestDelay               => ticd_CLK,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TO_X01((R_CLK_dly) AND (CE_ipd)) = '1',
          HeaderMsg               => InstancePath & "/DFFCR",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_CE_EQ_1_ANB_R_EQ_1_posedge or Tviol_CE_CLK_posedge or Tviol_R_CLK_CE_EQ_1_posedge or Pviol_CLK_CE_EQ_1_ANB_R_EQ_1;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => dffcetab,
        DataIn => (
               D_CLK_dly, CLK_dly,R_CLK_dly,'1', CE_CLK_dly));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (R_CLK_dly'last_event, tpd_R_Q, TRUE),
                 1 => (CLK_dly'last_event, tpd_CLK_Q, TRUE)),
       Mode => VitalInertial,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;

configuration CFG_DFFCR_VITAL of DFFCR is 
        for VITAL_VF
        end for; 
end CFG_DFFCR_VITAL;
----- VITAL model for cell DFFCRH -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;

LIBRARY VF1 ;
use VF1.VLOGTOVITAL_TABLES.all;



-- entity declaration --
entity DFFCRH is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_R_Q                        :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tsetup_D_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      thold_D_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      tsetup_CE_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      thold_CE_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      tpw_CLK_posedge 		:	VitalDelayType := 4.400 ns;
      tpw_R_posedge 		:	VitalDelayType := 4.400 ns;
      tperiod_CLK_posedge :	VitalDelayType := 8.800 ns;
      trecovery_R_CLK_negedge_posedge :	VitalDelayType := 2.200 ns;
      thold_R_CLK_negedge_posedge :	VitalDelayType := 2.200 ns;
      ticd_CLK                       :	VitalDelayType := 0.000 ns;
      tisd_D_CLK                     :	VitalDelayType := 0.000 ns;
      tisd_CE_CLK                     :	VitalDelayType := 0.000 ns;
      tisd_R_CLK                     :	VitalDelayType := 0.000 ns;
      tipd_CE                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_R                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      CE                             :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      R                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFFCRH : entity is TRUE;
end DFFCRH;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library VF1;
architecture VITAL_VF of DFFCRH is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL CE_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL R_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL D_CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL CE_CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL R_CLK_dly	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (CE_ipd, CE, tipd_CE);
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (R_ipd, R, tipd_R);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   VitalSignalDelay (CLK_dly, CLK_ipd, ticd_CLK);
   VitalSignalDelay (D_CLK_dly, D_ipd, tisd_D_CLK);
   VitalSignalDelay (CE_CLK_dly, CE_ipd, tisd_CE_CLK);
   VitalSignalDelay (R_CLK_dly, R_ipd, tisd_R_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (CE_ipd, CLK_dly, D_CLK_dly, R_CLK_dly, CE_CLK_dly)

   -- timing check results
   VARIABLE Tviol_D_CLK_CE_EQ_1_ANB_R_EQ_0_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_CE_EQ_1_ANB_R_EQ_0_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CE_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CE_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_R_CLK_CE_EQ_1_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_R_CLK_CE_EQ_1_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK_CE_EQ_1_ANB_R_EQ_0	: STD_ULOGIC := '0';
   VARIABLE Pviol_R				: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK_CE_EQ_1_ANB_R_EQ_0	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE PInfo_R				: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 4);
   VARIABLE R_inverted : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_CE_EQ_1_ANB_R_EQ_0_posedge,
          TimingData              => Tmkr_D_CLK_CE_EQ_1_ANB_R_EQ_0_posedge,
          TestSignal              => D_CLK_dly,
          TestSignalName          => "D",
          TestDelay               => tisd_D_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          SetupHigh               => tsetup_D_CLK_noedge_posedge,
          SetupLow                => tsetup_D_CLK_noedge_posedge,
          HoldHigh                => thold_D_CLK_noedge_posedge,
          HoldLow                 => thold_D_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(((NOT R_CLK_dly)) AND (CE_ipd)) = '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFFCRH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_CE_CLK_posedge,
          TimingData              => Tmkr_CE_CLK_posedge,
          TestSignal              => CE_CLK_dly,
          TestSignalName          => "CE",
          TestDelay               => tisd_CE_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          SetupHigh               => tsetup_CE_CLK_noedge_posedge,
          SetupLow                => tsetup_CE_CLK_noedge_posedge,
          HoldHigh                => thold_CE_CLK_noedge_posedge,
          HoldLow                 => thold_CE_CLK_noedge_posedge,
          CheckEnabled            => TRUE, 
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFFCRH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_R_CLK_CE_EQ_1_posedge,
          TimingData              => Tmkr_R_CLK_CE_EQ_1_posedge,
          TestSignal              => R_CLK_dly,
          TestSignalName          => "R",
          TestDelay               => tisd_R_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          Recovery                => trecovery_R_CLK_negedge_posedge,
          Removal                 => thold_R_CLK_negedge_posedge,
          ActiveLow               => FALSE,
          CheckEnabled            => 
                           TO_X01(CE_ipd) = '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFFCRH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_R,
          PeriodData              => PInfo_R,
          TestSignal              => R_CLK_dly,
          TestSignalName          => "R",
          TestDelay               => tisd_R_CLK,
          Period                  => 0 ns,
          PulseWidthHigh          => tpw_R_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => TRUE,
          HeaderMsg               => InstancePath & "/DFFCRH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK_CE_EQ_1_ANB_R_EQ_0,
          PeriodData              => PInfo_CLK_CE_EQ_1_ANB_R_EQ_0,
          TestSignal              => CLK_dly,
          TestSignalName          => "CLK",
          TestDelay               => ticd_CLK,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TO_X01(((NOT R_CLK_dly)) AND (CE_ipd)) = '1',
          HeaderMsg               => InstancePath & "/DFFCRH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_CE_EQ_1_ANB_R_EQ_0_posedge or Tviol_CE_CLK_posedge or Tviol_R_CLK_CE_EQ_1_posedge or Pviol_CLK_CE_EQ_1_ANB_R_EQ_0 or Pviol_R;
      R_inverted := (NOT R_CLK_dly);
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => dffcetab,
        DataIn => (
               D_CLK_dly, CLK_dly,R_inverted,'1', CE_CLK_dly));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (R_CLK_dly'last_event, tpd_R_Q, TRUE),
                 1 => (CLK_dly'last_event, tpd_CLK_Q, TRUE)),
       Mode => VitalInertial,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;

configuration CFG_DFFCRH_VITAL of DFFCRH is 
        for VITAL_VF
        end for; 
end CFG_DFFCRH_VITAL;
----- VITAL model for cell DFFCRS -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;

LIBRARY VF1 ;
use VF1.VLOGTOVITAL_TABLES.all;

-- entity declaration --
entity DFFCRS is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_S_Q                        :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tpd_R_Q                        :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tsetup_D_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      tsetup_CE_CLK_posedge_posedge :	VitalDelayType := 2.200 ns;
      thold_D_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      thold_CE_CLK_posedge_posedge :	VitalDelayType := 2.200 ns;
      tpw_CLK_posedge :	VitalDelayType := 4.400 ns;
      tperiod_CLK_posedge :	VitalDelayType := 8.800 ns;
      trecovery_R_CLK_posedge_posedge :	VitalDelayType := 2.200 ns;
      thold_R_CLK_posedge_posedge :	VitalDelayType := 2.200 ns;
      trecovery_S_CLK_posedge_posedge :	VitalDelayType := 2.200 ns;
      thold_S_CLK_posedge_posedge :	VitalDelayType := 2.200 ns;
      ticd_CLK                       :	VitalDelayType := 0.000 ns;
      tisd_D_CLK                     :	VitalDelayType := 0.000 ns;
      tisd_CE_CLK                     :	VitalDelayType := 0.000 ns;
      tisd_R_CLK                     :	VitalDelayType := 0.000 ns;
      tisd_S_CLK                     :	VitalDelayType := 0.000 ns;
      tipd_CE                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_R                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      CE                             :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      R                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFFCRS : entity is TRUE;
end DFFCRS;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library VF1;
architecture VITAL_VF of DFFCRS is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL CE_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL R_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL D_CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL R_CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL S_CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL CE_CLK_dly	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (CE_ipd, CE, tipd_CE);
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (R_ipd, R, tipd_R);
   VitalWireDelay (S_ipd, S, tipd_S);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   VitalSignalDelay (CLK_dly, CLK_ipd, ticd_CLK);
   VitalSignalDelay (D_CLK_dly, D_ipd, tisd_D_CLK);
   VitalSignalDelay (CE_CLK_dly, CE_ipd, tisd_CE_CLK);
   VitalSignalDelay (R_CLK_dly, R_ipd, tisd_R_CLK);
   VitalSignalDelay (S_CLK_dly, S_ipd, tisd_S_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (CE_CLK_dly, CLK_dly, D_CLK_dly, R_CLK_dly, S_CLK_dly)

   -- timing check results
   VARIABLE Tviol_D_CLK_CE_EQ_1_AN_R_EQ_1_AN_S_EQ_1_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_CE_EQ_1_AN_R_EQ_1_AN_S_EQ_1_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CE_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CE_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_R_CLK_CE_EQ_1_AN_S_EQ_1_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_R_CLK_CE_EQ_1_AN_S_EQ_1_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S_CLK_CE_EQ_1_AN_R_EQ_1_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S_CLK_CE_EQ_1_AN_R_EQ_1_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK_CE_EQ_1_AN_R_EQ_1_AN_S_EQ_1	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK_CE_EQ_1_AN_R_EQ_1_AN_S_EQ_1	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(1 to 5);
   VARIABLE CE_delayed : STD_ULOGIC := 'X';
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_CE_EQ_1_AN_R_EQ_1_AN_S_EQ_1_posedge,
          TimingData              => Tmkr_D_CLK_CE_EQ_1_AN_R_EQ_1_AN_S_EQ_1_posedge,
          TestSignal              => D_CLK_dly,
          TestSignalName          => "D",
          TestDelay               => tisd_D_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          SetupHigh               => tsetup_D_CLK_noedge_posedge,
          SetupLow                => tsetup_D_CLK_noedge_posedge,
          HoldHigh                => thold_D_CLK_noedge_posedge,
          HoldLow                 => thold_D_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((R_CLK_dly) AND (CE_CLK_dly) AND (S_CLK_dly))
                            /= '0',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFFCRS",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_CE_CLK_posedge,
          TimingData              => Tmkr_CE_CLK_posedge,
          TestSignal              => CE_CLK_dly,
          TestSignalName          => "CE",
          TestDelay               => tisd_CE_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          SetupHigh               => tsetup_CE_CLK_posedge_posedge,
          SetupLow                => tsetup_CE_CLK_posedge_posedge,
          HoldHigh                => thold_CE_CLK_posedge_posedge,
          HoldLow                 => thold_CE_CLK_posedge_posedge,
          CheckEnabled            => TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFFCRS",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_R_CLK_CE_EQ_1_AN_S_EQ_1_posedge,
          TimingData              => Tmkr_R_CLK_CE_EQ_1_AN_S_EQ_1_posedge,
          TestSignal              => R_CLK_dly,
          TestSignalName          => "R",
          TestDelay               => tisd_R_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          Recovery                => trecovery_R_CLK_posedge_posedge,
          Removal                 => thold_R_CLK_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TO_X01((S_CLK_dly) AND (CE_CLK_dly)) /= '0',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFFCRS",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_S_CLK_CE_EQ_1_AN_R_EQ_1_posedge,
          TimingData              => Tmkr_S_CLK_CE_EQ_1_AN_R_EQ_1_posedge,
          TestSignal              => S_CLK_dly,
          TestSignalName          => "S",
          TestDelay               => tisd_S_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          Recovery                => trecovery_S_CLK_posedge_posedge,
          Removal                 => thold_S_CLK_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TO_X01((R_CLK_dly) AND (CE_CLK_dly)) /= '0',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFFCRS",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK_CE_EQ_1_AN_R_EQ_1_AN_S_EQ_1,
          PeriodData              => PInfo_CLK_CE_EQ_1_AN_R_EQ_1_AN_S_EQ_1,
          TestSignal              => CLK_dly,
          TestSignalName          => "CLK",
          TestDelay               => ticd_CLK,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TO_X01(( (NOT S_CLK_dly) ) OR ( (NOT R_CLK_dly) )
                            ) /= '1',
          HeaderMsg               => InstancePath & "/DFFCRS",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_CE_EQ_1_AN_R_EQ_1_AN_S_EQ_1_posedge or Tviol_CE_CLK_posedge or Tviol_R_CLK_CE_EQ_1_AN_S_EQ_1_posedge or Pviol_CLK_CE_EQ_1_AN_R_EQ_1_AN_S_EQ_1 or Tviol_S_CLK_CE_EQ_1_AN_R_EQ_1_posedge;
      CE_delayed := CE_CLK_dly;
      D_delayed := D_CLK_dly;
      CLK_delayed := CLK_dly;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => dffcetab,
        DataIn => (
               D_delayed, CLK_delayed, R_CLK_dly, S_CLK_dly,CE_delayed ));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (S_CLK_dly'last_event, tpd_S_Q, TRUE),
                 1 => (R_CLK_dly'last_event, tpd_R_Q, TRUE),
                 2 => (CLK_dly'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;

configuration CFG_DFFCRS_VITAL of DFFCRS is 
        for VITAL_VF
        end for; 
end CFG_DFFCRS_VITAL;
----- VITAL model for cell DFFCRSH -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;
LIBRARY VF1 ;
use VF1.VLOGTOVITAL_TABLES.all;


-- entity declaration --
entity DFFCRSH is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_S_Q                        :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tpd_R_Q                        :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tsetup_D_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      thold_D_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      tsetup_CE_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      thold_CE_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      tpw_CLK_posedge :	VitalDelayType := 4.400 ns;
      tpw_R_posedge :	VitalDelayType := 4.400 ns;
      tpw_S_posedge :	VitalDelayType := 4.400 ns;
      tperiod_CLK_posedge :	VitalDelayType := 8.800 ns;
      trecovery_R_CLK_negedge_posedge :	VitalDelayType := 2.200 ns;
      thold_R_CLK_negedge_posedge :	VitalDelayType := 2.200 ns;
      trecovery_S_CLK_negedge_posedge :	VitalDelayType := 2.200 ns;
      thold_S_CLK_negedge_posedge :	VitalDelayType := 2.200 ns;
      ticd_CLK                       :	VitalDelayType := 0.000 ns;
      tisd_D_CLK                     :	VitalDelayType := 0.000 ns;
      tisd_R_CLK                     :	VitalDelayType := 0.000 ns;
      tisd_S_CLK                     :	VitalDelayType := 0.000 ns;
      tisd_CE_CLK                     :	VitalDelayType := 0.000 ns;
      tipd_CE                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_R                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      CE                             :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      R                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFFCRSH : entity is TRUE;
end DFFCRSH;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library VF1;
architecture VITAL_VF of DFFCRSH is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL CE_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL R_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL D_CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL R_CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL S_CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL CE_CLK_dly	 : STD_ULOGIC := 'X';


begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (CE_ipd, CE, tipd_CE);
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (R_ipd, R, tipd_R);
   VitalWireDelay (S_ipd, S, tipd_S);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   VitalSignalDelay (CLK_dly, CLK_ipd, ticd_CLK);
   VitalSignalDelay (D_CLK_dly, D_ipd, tisd_D_CLK);
   VitalSignalDelay (R_CLK_dly, R_ipd, tisd_R_CLK);
   VitalSignalDelay (S_CLK_dly, S_ipd, tisd_S_CLK);
   VitalSignalDelay (CE_CLK_dly, CE_ipd, tisd_CE_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (CE_CLK_dly, CLK_dly, D_CLK_dly, R_CLK_dly, S_CLK_dly)

   -- timing check results
   VARIABLE Tviol_D_CLK_CE_EQ_1_AN_R_EQ_0_AN_S_EQ_0_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_CE_EQ_1_AN_R_EQ_0_AN_S_EQ_0_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CE_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CE_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_R_CLK_CE_EQ_1_AN_S_EQ_0_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_R_CLK_CE_EQ_1_AN_S_EQ_0_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S_CLK_CE_EQ_1_AN_R_EQ_0_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S_CLK_CE_EQ_1_AN_R_EQ_0_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK_CE_EQ_1_AN_R_EQ_0_AN_S_EQ_0	: STD_ULOGIC := '0';
   VARIABLE Pviol_R	: STD_ULOGIC := '0';
   VARIABLE Pviol_S	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK_CE_EQ_1_AN_R_EQ_0_AN_S_EQ_0	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE PInfo_R	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE PInfo_S	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(1 to 5);
   VARIABLE CE_delayed : STD_ULOGIC := 'X';
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE R_inverted : STD_ULOGIC := 'X';
   VARIABLE S_inverted : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_CE_EQ_1_AN_R_EQ_0_AN_S_EQ_0_posedge,
          TimingData              => Tmkr_D_CLK_CE_EQ_1_AN_R_EQ_0_AN_S_EQ_0_posedge,
          TestSignal              => D_CLK_dly,
          TestSignalName          => "D",
          TestDelay               => tisd_D_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          SetupHigh               => tsetup_D_CLK_noedge_posedge,
          SetupLow                => tsetup_D_CLK_noedge_posedge,
          HoldHigh                => thold_D_CLK_noedge_posedge,
          HoldLow                 => thold_D_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(((NOT R_CLK_dly)) AND (CE_CLK_dly) AND ((NOT
                            S_CLK_dly))) /= '0',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFFCRSH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_CE_CLK_posedge,
          TimingData              => Tmkr_CE_CLK_posedge,
          TestSignal              => CE_CLK_dly,
          TestSignalName          => "CE",
          TestDelay               => tisd_CE_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          SetupHigh               => tsetup_CE_CLK_noedge_posedge,
          SetupLow                => tsetup_CE_CLK_noedge_posedge,
          HoldHigh                => thold_CE_CLK_noedge_posedge,
          HoldLow                 => thold_CE_CLK_noedge_posedge,
          CheckEnabled            => TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFFCRSH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_R_CLK_CE_EQ_1_AN_S_EQ_0_posedge,
          TimingData              => Tmkr_R_CLK_CE_EQ_1_AN_S_EQ_0_posedge,
          TestSignal              => R_CLK_dly,
          TestSignalName          => "R",
          TestDelay               => tisd_R_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          Recovery                => trecovery_R_CLK_negedge_posedge,
          Removal                 => thold_R_CLK_negedge_posedge,
          ActiveLow               => FALSE,
          CheckEnabled            => 
                           TO_X01(((NOT S_CLK_dly)) AND (CE_CLK_dly)) /= '0',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFFCRSH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_S_CLK_CE_EQ_1_AN_R_EQ_0_posedge,
          TimingData              => Tmkr_S_CLK_CE_EQ_1_AN_R_EQ_0_posedge,
          TestSignal              => S_CLK_dly,
          TestSignalName          => "S",
          TestDelay               => tisd_S_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          Recovery                => trecovery_S_CLK_negedge_posedge,
          Removal                 => thold_S_CLK_negedge_posedge,
          ActiveLow               => FALSE,
          CheckEnabled            => 
                           TO_X01(((NOT R_CLK_dly)) AND (CE_CLK_dly)) /= '0',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFFCRSH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_S,
          PeriodData              => PInfo_S,
          TestSignal              => S_CLK_dly,
          TestSignalName          => "S",
          TestDelay               => tisd_S_CLK,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_S_posedge,
          CheckEnabled            => TRUE, 
          HeaderMsg               => InstancePath & "/DFFCRSH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_R,
          PeriodData              => PInfo_R,
          TestSignal              => R_CLK_dly,
          TestSignalName          => "R",
          TestDelay               => tisd_R_CLK,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_R_posedge,
          CheckEnabled            => TRUE, 
          HeaderMsg               => InstancePath & "/DFFCRSH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK_CE_EQ_1_AN_R_EQ_0_AN_S_EQ_0,
          PeriodData              => PInfo_CLK_CE_EQ_1_AN_R_EQ_0_AN_S_EQ_0,
          TestSignal              => CLK_dly,
          TestSignalName          => "CLK",
          TestDelay               => ticd_CLK,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TO_X01(( S_CLK_dly ) OR ( R_CLK_dly ) ) /= '1',
          HeaderMsg               => InstancePath & "/DFFCRSH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_CE_EQ_1_AN_R_EQ_0_AN_S_EQ_0_posedge or Tviol_CE_CLK_posedge or Tviol_R_CLK_CE_EQ_1_AN_S_EQ_0_posedge or Tviol_S_CLK_CE_EQ_1_AN_R_EQ_0_posedge or Pviol_CLK_CE_EQ_1_AN_R_EQ_0_AN_S_EQ_0 or Pviol_R or Pviol_S;
      CE_delayed := CE_CLK_dly;
      D_delayed := D_CLK_dly;
      CLK_delayed := CLK_dly;
      R_inverted := (NOT R_CLK_dly);
      S_inverted := (NOT S_CLK_dly);
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => dffcetab,
        DataIn => (
               D_delayed, CLK_delayed,R_inverted,S_inverted,CE_delayed));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (S_CLK_dly'last_event, tpd_S_Q, TRUE),
                 1 => (R_CLK_dly'last_event, tpd_R_Q, TRUE),
                 2 => (CLK_dly'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;

configuration CFG_DFFCRSH_VITAL of DFFCRSH is 
        for VITAL_VF
        end for; 
end CFG_DFFCRSH_VITAL;
----- VITAL model for cell DFFCRSS -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;

LIBRARY VF1 ;
use VF1.VLOGTOVITAL_TABLES.all;



-- entity declaration --
entity DFFCRSS is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_S_Q                        :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tpd_R_Q                        :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tsetup_D_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      thold_D_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      tsetup_CE_CLK_posedge_posedge :	VitalDelayType := 2.200 ns;
      thold_CE_CLK_posedge_posedge :	VitalDelayType := 2.200 ns;
      tpw_CLK_posedge :	VitalDelayType := 4.400 ns;
      tperiod_CLK_posedge :	VitalDelayType := 8.800 ns;
      trecovery_R_CLK_posedge_posedge :	VitalDelayType := 2.200 ns;
      thold_R_CLK_posedge_posedge :	VitalDelayType := 2.200 ns;
      trecovery_S_CLK_posedge_posedge :	VitalDelayType := 2.200 ns;
      thold_S_CLK_posedge_posedge :	VitalDelayType := 2.200 ns;
      ticd_CLK                       :	VitalDelayType := 0.000 ns;
      tisd_D_CLK                     :	VitalDelayType := 0.000 ns;
      tisd_CE_CLK                     :	VitalDelayType := 0.000 ns;
      tisd_R_CLK                     :	VitalDelayType := 0.000 ns;
      tisd_S_CLK                     :	VitalDelayType := 0.000 ns;
      tipd_CE                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_R                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      CE                             :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      R                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFFCRSS : entity is TRUE;
end DFFCRSS;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library VF1;
architecture VITAL_VF of DFFCRSS is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL CE_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL R_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL D_CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL CE_CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL R_CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL S_CLK_dly	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (CE_ipd, CE, tipd_CE);
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (R_ipd, R, tipd_R);
   VitalWireDelay (S_ipd, S, tipd_S);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   VitalSignalDelay (CLK_dly, CLK_ipd, ticd_CLK);
   VitalSignalDelay (D_CLK_dly, D_ipd, tisd_D_CLK);
   VitalSignalDelay (CE_CLK_dly, CE_ipd, tisd_CE_CLK);
   VitalSignalDelay (R_CLK_dly, R_ipd, tisd_R_CLK);
   VitalSignalDelay (S_CLK_dly, S_ipd, tisd_S_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (CE_ipd, CLK_dly, D_CLK_dly, R_CLK_dly, S_CLK_dly, CE_CLK_dly)

   -- timing check results
   VARIABLE Tviol_D_CLK_CE_EQ_1_ANB_R_EQ_1_ANB_S_EQ_1_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_CE_EQ_1_ANB_R_EQ_1_ANB_S_EQ_1_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CE_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CE_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_R_CLK_CE_EQ_1_ANB_S_EQ_1_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_R_CLK_CE_EQ_1_ANB_S_EQ_1_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S_CLK_CE_EQ_1_ANB_R_EQ_1_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S_CLK_CE_EQ_1_ANB_R_EQ_1_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK_CE_EQ_1_ANB_R_EQ_1_ANB_S_EQ_1	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK_CE_EQ_1_ANB_R_EQ_1_ANB_S_EQ_1	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE D_int : STD_ULOGIC ;
   VARIABLE S_inverted : STD_ULOGIC ;
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 4);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_CE_EQ_1_ANB_R_EQ_1_ANB_S_EQ_1_posedge,
          TimingData              => Tmkr_D_CLK_CE_EQ_1_ANB_R_EQ_1_ANB_S_EQ_1_posedge,
          TestSignal              => D_CLK_dly,
          TestSignalName          => "D",
          TestDelay               => tisd_D_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          SetupHigh               => tsetup_D_CLK_noedge_posedge,
          SetupLow                => tsetup_D_CLK_noedge_posedge,
          HoldHigh                => thold_D_CLK_noedge_posedge,
          HoldLow                 => thold_D_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((R_CLK_dly) AND (CE_ipd) AND (S_CLK_dly)) = '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFFCRSS",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_CE_CLK_posedge,
          TimingData              => Tmkr_CE_CLK_posedge,
          TestSignal              => CE_CLK_dly,
          TestSignalName          => "CE",
          TestDelay               => tisd_CE_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          SetupHigh               => tsetup_CE_CLK_posedge_posedge,
          SetupLow                => tsetup_CE_CLK_posedge_posedge,
          HoldHigh                => thold_CE_CLK_posedge_posedge,
          HoldLow                 => thold_CE_CLK_posedge_posedge,
          CheckEnabled            => TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFFCRSS",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_R_CLK_CE_EQ_1_ANB_S_EQ_1_posedge,
          TimingData              => Tmkr_R_CLK_CE_EQ_1_ANB_S_EQ_1_posedge,
          TestSignal              => R_CLK_dly,
          TestSignalName          => "R",
          TestDelay               => tisd_R_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          Recovery                => trecovery_R_CLK_posedge_posedge,
          Removal                 => thold_R_CLK_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TO_X01((S_CLK_dly) AND (CE_ipd)) = '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFFCRSS",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_S_CLK_CE_EQ_1_ANB_R_EQ_1_posedge,
          TimingData              => Tmkr_S_CLK_CE_EQ_1_ANB_R_EQ_1_posedge,
          TestSignal              => S_CLK_dly,
          TestSignalName          => "S",
          TestDelay               => tisd_S_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          Recovery                => trecovery_S_CLK_posedge_posedge,
          Removal                 => thold_S_CLK_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TO_X01((R_CLK_dly) AND (CE_ipd)) = '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFFCRSS",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK_CE_EQ_1_ANB_R_EQ_1_ANB_S_EQ_1,
          PeriodData              => PInfo_CLK_CE_EQ_1_ANB_R_EQ_1_ANB_S_EQ_1,
          TestSignal              => CLK_dly,
          TestSignalName          => "CLK",
          TestDelay               => ticd_CLK,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TO_X01((R_CLK_dly) AND (CE_ipd) AND (S_CLK_dly)) = '1',
          HeaderMsg               => InstancePath & "/DFFCRSS",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_CE_EQ_1_ANB_R_EQ_1_ANB_S_EQ_1_posedge or Tviol_CE_CLK_posedge or Tviol_R_CLK_CE_EQ_1_ANB_S_EQ_1_posedge or Tviol_S_CLK_CE_EQ_1_ANB_R_EQ_1_posedge or Pviol_CLK_CE_EQ_1_ANB_R_EQ_1_ANB_S_EQ_1;
      S_inverted := VitalINV (S_CLK_dly);
      D_int := VitalOR2 (D_CLK_dly,S_inverted);
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => dffcetab,
        DataIn => (
               D_int, CLK_dly, R_CLK_dly, '1', CE_CLK_dly));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (S_CLK_dly'last_event, tpd_S_Q, TRUE),
                 1 => (R_CLK_dly'last_event, tpd_R_Q, TRUE),
                 2 => (CLK_dly'last_event, tpd_CLK_Q, TRUE)),
       Mode => VitalInertial,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;

configuration CFG_DFFCRSS_VITAL of DFFCRSS is 
        for VITAL_VF
        end for; 
end CFG_DFFCRSS_VITAL;
----- VITAL model for cell DFFCRSSH -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;

LIBRARY VF1 ;
use VF1.VLOGTOVITAL_TABLES.all;



-- entity declaration --
entity DFFCRSSH is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_S_Q                        :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tpd_R_Q                        :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tsetup_D_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      thold_D_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      tsetup_CE_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      thold_CE_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      tpw_CLK_posedge :	VitalDelayType := 4.400 ns;
      tpw_R_posedge :	VitalDelayType := 4.400 ns;
      tperiod_CLK_posedge :	VitalDelayType := 8.800 ns;
      trecovery_R_CLK_negedge_posedge :	VitalDelayType := 2.200 ns;
      thold_R_CLK_negedge_posedge :	VitalDelayType := 2.200 ns;
      tsetup_S_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      thold_S_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      ticd_CLK                       :	VitalDelayType := 0.000 ns;
      tisd_D_CLK                     :	VitalDelayType := 0.000 ns;
      tisd_CE_CLK                     :	VitalDelayType := 0.000 ns;
      tisd_R_CLK                     :	VitalDelayType := 0.000 ns;
      tisd_S_CLK                     :	VitalDelayType := 0.000 ns;
      tipd_CE                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_R                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      CE                             :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      R                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFFCRSSH : entity is TRUE;
end DFFCRSSH;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library VF1;
architecture VITAL_VF of DFFCRSSH is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL CE_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL R_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL D_CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL CE_CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL R_CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL S_CLK_dly	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (CE_ipd, CE, tipd_CE);
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (R_ipd, R, tipd_R);
   VitalWireDelay (S_ipd, S, tipd_S);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   VitalSignalDelay (CLK_dly, CLK_ipd, ticd_CLK);
   VitalSignalDelay (D_CLK_dly, D_ipd, tisd_D_CLK);
   VitalSignalDelay (CE_CLK_dly, CE_ipd, tisd_CE_CLK);
   VitalSignalDelay (R_CLK_dly, R_ipd, tisd_R_CLK);
   VitalSignalDelay (S_CLK_dly, S_ipd, tisd_S_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (CE_ipd, CLK_dly, D_CLK_dly, R_CLK_dly, S_CLK_dly, CE_CLK_dly)

   -- timing check results
   VARIABLE Tviol_D_CLK_CE_EQ_1_ANB_R_EQ_0_ANB_S_EQ_0_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_CE_EQ_1_ANB_R_EQ_0_ANB_S_EQ_0_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CE_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CE_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_R_CLK_CE_EQ_1_ANB_S_EQ_0_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_R_CLK_CE_EQ_1_ANB_S_EQ_0_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S_CLK_CE_EQ_1_ANB_R_EQ_0_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S_CLK_CE_EQ_1_ANB_R_EQ_0_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK_CE_EQ_1_ANB_R_EQ_0_ANB_S_EQ_0	: STD_ULOGIC := '0';
   VARIABLE Pviol_R	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK_CE_EQ_1_ANB_R_EQ_0_ANB_S_EQ_0	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE PInfo_R	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 4);
   VARIABLE R_inverted : STD_ULOGIC := 'X';
   VARIABLE D_int : STD_ULOGIC := '0';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_CE_EQ_1_ANB_R_EQ_0_ANB_S_EQ_0_posedge,
          TimingData              => Tmkr_D_CLK_CE_EQ_1_ANB_R_EQ_0_ANB_S_EQ_0_posedge,
          TestSignal              => D_CLK_dly,
          TestSignalName          => "D",
          TestDelay               => tisd_D_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          SetupHigh               => tsetup_D_CLK_noedge_posedge,
          SetupLow                => tsetup_D_CLK_noedge_posedge,
          HoldHigh                => thold_D_CLK_noedge_posedge,
          HoldLow                 => thold_D_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(((NOT R_CLK_dly)) AND (CE_ipd) AND ((NOT S_CLK_dly))) = '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFFCRSSH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_CE_CLK_posedge,
          TimingData              => Tmkr_CE_CLK_posedge,
          TestSignal              => CE_CLK_dly,
          TestSignalName          => "CE",
          TestDelay               => tisd_CE_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          SetupHigh               => tsetup_CE_CLK_noedge_posedge,
          SetupLow                => tsetup_CE_CLK_noedge_posedge,
          HoldHigh                => thold_CE_CLK_noedge_posedge,
          HoldLow                 => thold_CE_CLK_noedge_posedge,
          CheckEnabled            => TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFFCRSSH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_R_CLK_CE_EQ_1_ANB_S_EQ_0_posedge,
          TimingData              => Tmkr_R_CLK_CE_EQ_1_ANB_S_EQ_0_posedge,
          TestSignal              => R_CLK_dly,
          TestSignalName          => "R",
          TestDelay               => tisd_R_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          Recovery                => trecovery_R_CLK_negedge_posedge,
          Removal                 => thold_R_CLK_negedge_posedge,
          ActiveLow               => FALSE,
          CheckEnabled            => 
                           TO_X01(((NOT S_CLK_dly)) AND (CE_ipd)) = '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFFCRSSH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_S_CLK_CE_EQ_1_ANB_R_EQ_0_posedge,
          TimingData              => Tmkr_S_CLK_CE_EQ_1_ANB_R_EQ_0_posedge,
          TestSignal              => S_CLK_dly,
          TestSignalName          => "S",
          TestDelay               => tisd_S_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          SetupHigh               => tsetup_S_CLK_noedge_posedge,
          SetupLow                => tsetup_S_CLK_noedge_posedge,
          HoldHigh                => thold_S_CLK_noedge_posedge,
          HoldLow                 => thold_S_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(((NOT R_CLK_dly)) AND (CE_ipd)) = '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFFCRSSH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_R,
          PeriodData              => PInfo_R,
          TestSignal              => R_CLK_dly,
          TestSignalName          => "R",
          TestDelay               => tisd_R_CLK,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_R_posedge,
          CheckEnabled            => TRUE, 
          HeaderMsg               => InstancePath & "/DFFCRSSH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK_CE_EQ_1_ANB_R_EQ_0_ANB_S_EQ_0,
          PeriodData              => PInfo_CLK_CE_EQ_1_ANB_R_EQ_0_ANB_S_EQ_0,
          TestSignal              => CLK_dly,
          TestSignalName          => "CLK",
          TestDelay               => ticd_CLK,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TO_X01(((NOT R_CLK_dly)) AND (CE_ipd) AND ((NOT S_CLK_dly))) = '1',
          HeaderMsg               => InstancePath & "/DFFCRSSH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_CE_EQ_1_ANB_R_EQ_0_ANB_S_EQ_0_posedge or Tviol_CE_CLK_posedge or Tviol_R_CLK_CE_EQ_1_ANB_S_EQ_0_posedge or Tviol_S_CLK_CE_EQ_1_ANB_R_EQ_0_posedge or Pviol_CLK_CE_EQ_1_ANB_R_EQ_0_ANB_S_EQ_0 or Pviol_R;
      R_inverted := (NOT R_CLK_dly);
      D_int := VitalOR2 (D_CLK_dly,S_CLK_dly);
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => dffcetab,
        DataIn => (
               D_int, CLK_dly, R_inverted, '1', CE_CLK_dly));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (S_CLK_dly'last_event, tpd_S_Q, TRUE),
                 1 => (R_CLK_dly'last_event, tpd_R_Q, TRUE),
                 2 => (CLK_dly'last_event, tpd_CLK_Q, TRUE)),
       Mode => VitalInertial,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;

configuration CFG_DFFCRSSH_VITAL of DFFCRSSH is 
        for VITAL_VF
        end for; 
end CFG_DFFCRSSH_VITAL;
----- VITAL model for cell DFFCS -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;

LIBRARY VF1 ;
use VF1.VLOGTOVITAL_TABLES.all;



-- entity declaration --
entity DFFCS is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_S_Q                        :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tsetup_D_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      thold_D_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      tsetup_CE_CLK_posedge_posedge :	VitalDelayType := 2.200 ns;
      thold_CE_CLK_posedge_posedge :	VitalDelayType := 2.200 ns;
      tpw_CLK_posedge :	VitalDelayType := 4.400 ns;
      tperiod_CLK_posedge :	VitalDelayType := 8.800 ns;
      trecovery_S_CLK_posedge_posedge :	VitalDelayType := 2.200 ns;
      thold_S_CLK_posedge_posedge :	VitalDelayType := 2.200 ns;
      ticd_CLK                       :	VitalDelayType := 0.000 ns;
      tisd_D_CLK                     :	VitalDelayType := 0.000 ns;
      tisd_CE_CLK                     :	VitalDelayType := 0.000 ns;
      tisd_S_CLK                     :	VitalDelayType := 0.000 ns;
      tipd_CE                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      CE                             :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFFCS : entity is TRUE;
end DFFCS;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library VF1;
architecture VITAL_VF of DFFCS is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL CE_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL D_CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL CE_CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL S_CLK_dly	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (CE_ipd, CE, tipd_CE);
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (S_ipd, S, tipd_S);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   VitalSignalDelay (CLK_dly, CLK_ipd, ticd_CLK);
   VitalSignalDelay (D_CLK_dly, D_ipd, tisd_D_CLK);
   VitalSignalDelay (CE_CLK_dly, CE_ipd, tisd_CE_CLK);
   VitalSignalDelay (S_CLK_dly, S_ipd, tisd_S_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (CE_ipd, CLK_dly, D_CLK_dly, S_CLK_dly, CE_CLK_dly)

   -- timing check results
   VARIABLE Tviol_D_CLK_CE_EQ_1_ANB_S_EQ_1_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_CE_EQ_1_ANB_S_EQ_1_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CE_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CE_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S_CLK_CE_EQ_1_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S_CLK_CE_EQ_1_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK_CE_EQ_1_ANB_S_EQ_1	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK_CE_EQ_1_ANB_S_EQ_1	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 4);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_CE_EQ_1_ANB_S_EQ_1_posedge,
          TimingData              => Tmkr_D_CLK_CE_EQ_1_ANB_S_EQ_1_posedge,
          TestSignal              => D_CLK_dly,
          TestSignalName          => "D",
          TestDelay               => tisd_D_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          SetupHigh               => tsetup_D_CLK_noedge_posedge,
          SetupLow                => tsetup_D_CLK_noedge_posedge,
          HoldHigh                => thold_D_CLK_noedge_posedge,
          HoldLow                 => thold_D_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((S_CLK_dly) AND (CE_ipd)) = '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFFCS",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_CE_CLK_posedge,
          TimingData              => Tmkr_CE_CLK_posedge,
          TestSignal              => CE_CLK_dly,
          TestSignalName          => "CE",
          TestDelay               => tisd_CE_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          SetupHigh               => tsetup_CE_CLK_posedge_posedge,
          SetupLow                => tsetup_CE_CLK_posedge_posedge,
          HoldHigh                => thold_CE_CLK_posedge_posedge,
          HoldLow                 => thold_CE_CLK_posedge_posedge,
          CheckEnabled            => TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFFCS",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_S_CLK_CE_EQ_1_posedge,
          TimingData              => Tmkr_S_CLK_CE_EQ_1_posedge,
          TestSignal              => S_CLK_dly,
          TestSignalName          => "S",
          TestDelay               => tisd_S_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          Recovery                => trecovery_S_CLK_posedge_posedge,
          Removal                 => thold_S_CLK_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TO_X01(CE_ipd) = '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFFCS",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK_CE_EQ_1_ANB_S_EQ_1,
          PeriodData              => PInfo_CLK_CE_EQ_1_ANB_S_EQ_1,
          TestSignal              => CLK_dly,
          TestSignalName          => "CLK",
          TestDelay               => ticd_CLK,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                          TO_X01((S_CLK_dly) AND (CE_ipd)) = '1',
          HeaderMsg               => InstancePath & "/DFFCS",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_CE_EQ_1_ANB_S_EQ_1_posedge or Tviol_CE_CLK_posedge or Tviol_S_CLK_CE_EQ_1_posedge or Pviol_CLK_CE_EQ_1_ANB_S_EQ_1;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => dffcetab,
        DataIn => (
               D_CLK_dly, CLK_dly,'1',S_CLK_dly, CE_CLK_dly));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (S_CLK_dly'last_event, tpd_S_Q, TRUE),
                 1 => (CLK_dly'last_event, tpd_CLK_Q, TRUE)),
       Mode => VitalInertial,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;

configuration CFG_DFFCS_VITAL of DFFCS is 
        for VITAL_VF
        end for; 
end CFG_DFFCS_VITAL;
----- VITAL model for cell DFFCSH -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;

LIBRARY VF1 ;
use VF1.VLOGTOVITAL_TABLES.all;



-- entity declaration --
entity DFFCSH is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_S_Q                        :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tsetup_D_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      thold_D_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      tsetup_CE_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      thold_CE_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      tpw_CLK_posedge :	VitalDelayType := 4.400 ns;
      tpw_S_posedge :	VitalDelayType := 4.400 ns;
      tperiod_CLK_posedge :	VitalDelayType := 8.800 ns;
      trecovery_S_CLK_negedge_posedge :	VitalDelayType := 2.200 ns;
      thold_S_CLK_negedge_posedge :	VitalDelayType := 2.200 ns;
      ticd_CLK                       :	VitalDelayType := 0.000 ns;
      tisd_D_CLK                     :	VitalDelayType := 0.000 ns;
      tisd_CE_CLK                     :	VitalDelayType := 0.000 ns;
      tisd_S_CLK                     :	VitalDelayType := 0.000 ns;
      tipd_CE                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      CE                             :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFFCSH : entity is TRUE;
end DFFCSH;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library VF1;
architecture VITAL_VF of DFFCSH is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL CE_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL D_CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL CE_CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL S_CLK_dly	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (CE_ipd, CE, tipd_CE);
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (S_ipd, S, tipd_S);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   VitalSignalDelay (CLK_dly, CLK_ipd, ticd_CLK);
   VitalSignalDelay (D_CLK_dly, D_ipd, tisd_D_CLK);
   VitalSignalDelay (CE_CLK_dly, CE_ipd, tisd_CE_CLK);
   VitalSignalDelay (S_CLK_dly, S_ipd, tisd_S_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (CE_ipd, CLK_dly, D_CLK_dly, S_CLK_dly, CE_CLK_dly)

   -- timing check results
   VARIABLE Tviol_D_CLK_CE_EQ_1_ANB_S_EQ_0_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_CE_EQ_1_ANB_S_EQ_0_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CE_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CE_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S_CLK_CE_EQ_1_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S_CLK_CE_EQ_1_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK_CE_EQ_1_ANB_S_EQ_0	: STD_ULOGIC := '0';
   VARIABLE Pviol_S	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK_CE_EQ_1_ANB_S_EQ_0	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE PInfo_S	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 4);
   VARIABLE S_inverted : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_CE_EQ_1_ANB_S_EQ_0_posedge,
          TimingData              => Tmkr_D_CLK_CE_EQ_1_ANB_S_EQ_0_posedge,
          TestSignal              => D_CLK_dly,
          TestSignalName          => "D",
          TestDelay               => tisd_D_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          SetupHigh               => tsetup_D_CLK_noedge_posedge,
          SetupLow                => tsetup_D_CLK_noedge_posedge,
          HoldHigh                => thold_D_CLK_noedge_posedge,
          HoldLow                 => thold_D_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(((NOT S_CLK_dly)) AND (CE_ipd)) = '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFFCSH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_CE_CLK_posedge,
          TimingData              => Tmkr_CE_CLK_posedge,
          TestSignal              => CE_CLK_dly,
          TestSignalName          => "CE",
          TestDelay               => tisd_CE_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          SetupHigh               => tsetup_CE_CLK_noedge_posedge,
          SetupLow                => tsetup_CE_CLK_noedge_posedge,
          HoldHigh                => thold_CE_CLK_noedge_posedge,
          HoldLow                 => thold_CE_CLK_noedge_posedge,
          CheckEnabled            => TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFFCSH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_S_CLK_CE_EQ_1_posedge,
          TimingData              => Tmkr_S_CLK_CE_EQ_1_posedge,
          TestSignal              => S_CLK_dly,
          TestSignalName          => "S",
          TestDelay               => tisd_S_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          Recovery                => trecovery_S_CLK_negedge_posedge,
          Removal                 => thold_S_CLK_negedge_posedge,
          ActiveLow               => FALSE,
          CheckEnabled            => 
                           TO_X01(CE_ipd) = '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFFCSH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_S,
          PeriodData              => PInfo_S,
          TestSignal              => S_CLK_dly,
          TestSignalName          => "S",
          TestDelay               => tisd_S_CLK,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_S_posedge,
          CheckEnabled            => TRUE, 
          HeaderMsg               => InstancePath & "/DFFCSH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK_CE_EQ_1_ANB_S_EQ_0,
          PeriodData              => PInfo_CLK_CE_EQ_1_ANB_S_EQ_0,
          TestSignal              => CLK_dly,
          TestSignalName          => "CLK",
          TestDelay               => ticd_CLK,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TO_X01(((NOT S_CLK_dly)) AND (CE_ipd)) = '1',
          HeaderMsg               => InstancePath & "/DFFCSH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_CE_EQ_1_ANB_S_EQ_0_posedge or Tviol_CE_CLK_posedge or Tviol_S_CLK_CE_EQ_1_posedge or Pviol_CLK_CE_EQ_1_ANB_S_EQ_0 or Pviol_S;
      S_inverted := (NOT S_CLK_dly);
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => dffcetab,
        DataIn => (
               D_CLK_dly, CLK_dly,'1', S_inverted, CE_CLK_dly));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (S_CLK_dly'last_event, tpd_S_Q, TRUE),
                 1 => (CLK_dly'last_event, tpd_CLK_Q, TRUE)),
       Mode => VitalInertial,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;

configuration CFG_DFFCSH_VITAL of DFFCSH is 
        for VITAL_VF
        end for; 
end CFG_DFFCSH_VITAL;
----- VITAL model for cell DFFR -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;

LIBRARY VF1 ;
use VF1.VLOGTOVITAL_TABLES.all;



-- entity declaration --
entity DFFR is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_R_Q                        :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tsetup_D_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      thold_D_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      tpw_CLK_posedge         :	VitalDelayType := 4.400 ns;
      tperiod_CLK_posedge             :	VitalDelayType := 8.800 ns;
      trecovery_R_CLK_posedge_posedge :	VitalDelayType := 2.200 ns;
      thold_R_CLK_posedge_posedge    :	VitalDelayType := 2.200 ns;
      ticd_CLK                       :	VitalDelayType := 0.000 ns;
      tisd_D_CLK                     :	VitalDelayType := 0.000 ns;
      tisd_R_CLK                     :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_R                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      R                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFFR : entity is TRUE;
end DFFR;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library VF1;
architecture VITAL_VF of DFFR is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL R_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL D_CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL R_CLK_dly	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (R_ipd, R, tipd_R);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   VitalSignalDelay (CLK_dly, CLK_ipd, ticd_CLK);
   VitalSignalDelay (D_CLK_dly, D_ipd, tisd_D_CLK);
   VitalSignalDelay (R_CLK_dly, R_ipd, tisd_R_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (CLK_dly, D_CLK_dly, R_CLK_dly)

   -- timing check results
   VARIABLE Tviol_D_CLK_R_EQ_1_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_R_EQ_1_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_R_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_R_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK_R_EQ_1	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK_R_EQ_1	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 3);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_R_EQ_1_posedge,
          TimingData              => Tmkr_D_CLK_R_EQ_1_posedge,
          TestSignal              => D_CLK_dly,
          TestSignalName          => "D",
          TestDelay               => tisd_D_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          SetupHigh               => tsetup_D_CLK_noedge_posedge,
          SetupLow                => tsetup_D_CLK_noedge_posedge,
          HoldHigh                => thold_D_CLK_noedge_posedge,
          HoldLow                 => thold_D_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(R_CLK_dly) = '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFFR",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_R_CLK_posedge,
          TimingData              => Tmkr_R_CLK_posedge,
          TestSignal              => R_CLK_dly,
          TestSignalName          => "R",
          TestDelay               => tisd_R_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          Recovery                => trecovery_R_CLK_posedge_posedge,
          Removal                 => thold_R_CLK_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFFR",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK_R_EQ_1,
          PeriodData              => PInfo_CLK_R_EQ_1,
          TestSignal              => CLK_dly,
          TestSignalName          => "CLK",
          TestDelay               => ticd_CLK,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TO_X01((R_CLK_dly) ) = '1',
          HeaderMsg               => InstancePath & "/DFFR",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_R_EQ_1_posedge or Tviol_R_CLK_posedge or Pviol_CLK_R_EQ_1;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => dfftab,
        DataIn => (
              D_CLK_dly, CLK_dly, R_CLK_dly, '1'));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (R_CLK_dly'last_event, tpd_R_Q, TRUE),
                 1 => (CLK_dly'last_event, tpd_CLK_Q, TRUE)),
       Mode => VitalInertial,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;

configuration CFG_DFFR_VITAL of DFFR is 
        for VITAL_VF
        end for; 
end CFG_DFFR_VITAL;
----- VITAL model for cell DFFRH -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;

LIBRARY VF1 ;
use VF1.VLOGTOVITAL_TABLES.all;



-- entity declaration --
entity DFFRH is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_R_Q                        :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tsetup_D_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      thold_D_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      tpw_CLK_posedge         :	VitalDelayType := 4.400 ns;
      tpw_R_posedge         :	VitalDelayType := 4.400 ns;
      tperiod_CLK_posedge             :	VitalDelayType := 8.800 ns;
      trecovery_R_CLK_negedge_posedge :	VitalDelayType := 2.200 ns;
      thold_R_CLK_negedge_posedge    :	VitalDelayType := 2.200 ns;
      ticd_CLK                       :	VitalDelayType := 0.000 ns;
      tisd_D_CLK                     :	VitalDelayType := 0.000 ns;
      tisd_R_CLK                     :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_R                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      R                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFFRH : entity is TRUE;
end DFFRH;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library VF1;
architecture VITAL_VF of DFFRH is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL R_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL D_CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL R_CLK_dly	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (R_ipd, R, tipd_R);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   VitalSignalDelay (CLK_dly, CLK_ipd, ticd_CLK);
   VitalSignalDelay (D_CLK_dly, D_ipd, tisd_D_CLK);
   VitalSignalDelay (R_CLK_dly, R_ipd, tisd_R_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (CLK_dly, D_CLK_dly, R_CLK_dly)

   -- timing check results
   VARIABLE Tviol_D_CLK_R_EQ_0_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_R_EQ_0_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_R_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_R_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK_R_EQ_0	: STD_ULOGIC := '0';
   VARIABLE Pviol_R	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK_R_EQ_0	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE PInfo_R	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 3);
   VARIABLE R_inverted : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_R_EQ_0_posedge,
          TimingData              => Tmkr_D_CLK_R_EQ_0_posedge,
          TestSignal              => D_CLK_dly,
          TestSignalName          => "D",
          TestDelay               => tisd_D_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          SetupHigh               => tsetup_D_CLK_noedge_posedge,
          SetupLow                => tsetup_D_CLK_noedge_posedge,
          HoldHigh                => thold_D_CLK_noedge_posedge,
          HoldLow                 => thold_D_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((R_CLK_dly)) = '0',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFFRH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_R_CLK_posedge,
          TimingData              => Tmkr_R_CLK_posedge,
          TestSignal              => R_CLK_dly,
          TestSignalName          => "R",
          TestDelay               => tisd_R_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          Recovery                => trecovery_R_CLK_negedge_posedge,
          Removal                 => thold_R_CLK_negedge_posedge,
          ActiveLow               => FALSE,
          CheckEnabled            => TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFFRH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_R,
          PeriodData              => PInfo_R,
          TestSignal              => R_CLK_dly,
          TestSignalName          => "R",
          TestDelay               => tisd_R_CLK,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_R_posedge,
          CheckEnabled            => TRUE, 
          HeaderMsg               => InstancePath & "/DFFRH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK_R_EQ_0,
          PeriodData              => PInfo_CLK_R_EQ_0,
          TestSignal              => CLK_dly,
          TestSignalName          => "CLK",
          TestDelay               => ticd_CLK,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TO_X01(R_CLK_dly ) = '0',
          HeaderMsg               => InstancePath & "/DFFRH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_R_EQ_0_posedge or Tviol_R_CLK_posedge or Pviol_CLK_R_EQ_0 or Pviol_R;
      R_inverted := (NOT R_CLK_dly);
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => dfftab,
        DataIn => (
               D_CLK_dly, CLK_dly, R_inverted, '1'));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (R_CLK_dly'last_event, tpd_R_Q, TRUE),
                 1 => (CLK_dly'last_event, tpd_CLK_Q, TRUE)),
       Mode => VitalInertial,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;

configuration CFG_DFFRH_VITAL of DFFRH is 
        for VITAL_VF
        end for; 
end CFG_DFFRH_VITAL;
----- VITAL model for cell DFFRS -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;
LIBRARY VF1 ;
use VF1.VLOGTOVITAL_TABLES.all;

-- entity declaration --
entity DFFRS is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_R_Q                        :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tpd_S_Q                        :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tsetup_D_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      thold_D_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      tpw_CLK_posedge :	VitalDelayType := 4.400 ns;
      tpw_R_negedge :	VitalDelayType := 4.400 ns;
      tpw_S_negedge :	VitalDelayType := 4.400 ns;
      tperiod_CLK_posedge   :	VitalDelayType := 8.800 ns;
      trecovery_R_CLK_posedge_posedge :	VitalDelayType := 2.200 ns;
      thold_R_CLK_posedge_posedge :	VitalDelayType := 2.200 ns;
      trecovery_S_CLK_posedge_posedge :	VitalDelayType := 2.200 ns;
      thold_S_CLK_posedge_posedge :	VitalDelayType := 2.200 ns;
      ticd_CLK                       :	VitalDelayType := 0.000 ns;
      tisd_D_CLK                     :	VitalDelayType := 0.000 ns;
      tisd_R_CLK                     :	VitalDelayType := 0.000 ns;
      tisd_S_CLK                     :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_R                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      R                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFFRS : entity is TRUE;
end DFFRS;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library VF1;
architecture VITAL_VF of DFFRS is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL R_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL D_CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL R_CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL S_CLK_dly	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (R_ipd, R, tipd_R);
   VitalWireDelay (S_ipd, S, tipd_S);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   VitalSignalDelay (CLK_dly, CLK_ipd, ticd_CLK);
   VitalSignalDelay (D_CLK_dly, D_ipd, tisd_D_CLK);
   VitalSignalDelay (R_CLK_dly, R_ipd, tisd_R_CLK);
   VitalSignalDelay (S_CLK_dly, S_ipd, tisd_S_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (CLK_dly, D_CLK_dly, R_CLK_dly, S_CLK_dly)

   -- timing check results
   VARIABLE Tviol_D_CLK_R_EQ_1_AN_S_EQ_1_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_R_EQ_1_AN_S_EQ_1_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_R_CLK_S_EQ_1_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_R_CLK_S_EQ_1_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S_CLK_R_EQ_1_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S_CLK_R_EQ_1_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK_R_EQ_1_AN_S_EQ_1	: STD_ULOGIC := '0';
   VARIABLE Pviol_R			: STD_ULOGIC := '0';
   VARIABLE Pviol_S			: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK_R_EQ_1_AN_S_EQ_1	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE PInfo_R			: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE PInfo_S			: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(1 to 4);
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_R_EQ_1_AN_S_EQ_1_posedge,
          TimingData              => Tmkr_D_CLK_R_EQ_1_AN_S_EQ_1_posedge,
          TestSignal              => D_CLK_dly,
          TestSignalName          => "D",
          TestDelay               => tisd_D_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          SetupHigh               => tsetup_D_CLK_noedge_posedge,
          SetupLow                => tsetup_D_CLK_noedge_posedge,
          HoldHigh                => thold_D_CLK_noedge_posedge,
          HoldLow                 => thold_D_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((S_CLK_dly) AND (R_CLK_dly)) /= '0',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFFRS",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_R_CLK_S_EQ_1_posedge,
          TimingData              => Tmkr_R_CLK_S_EQ_1_posedge,
          TestSignal              => R_CLK_dly,
          TestSignalName          => "R",
          TestDelay               => tisd_R_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          Recovery                => trecovery_R_CLK_posedge_posedge,
          Removal                 => thold_R_CLK_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TO_X01(S_CLK_dly) /= '0',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFFRS",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_S_CLK_R_EQ_1_posedge,
          TimingData              => Tmkr_S_CLK_R_EQ_1_posedge,
          TestSignal              => S_CLK_dly,
          TestSignalName          => "S",
          TestDelay               => tisd_S_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          Recovery                => trecovery_S_CLK_posedge_posedge,
          Removal                 => thold_S_CLK_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TO_X01(R_CLK_dly) /= '0',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFFRS",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_S,
          PeriodData              => PInfo_S,
          TestSignal              => S_CLK_dly,
          TestSignalName          => "S",
          TestDelay               => tisd_S_CLK,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_S_negedge,
          CheckEnabled            => TRUE,
          HeaderMsg               => InstancePath & "/DFFRS",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_R,
          PeriodData              => PInfo_R,
          TestSignal              => R_CLK_dly,
          TestSignalName          => "R",
          TestDelay               => tisd_R_CLK,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_R_negedge,
          CheckEnabled            => TRUE, 
          HeaderMsg               => InstancePath & "/DFFRS",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK_R_EQ_1_AN_S_EQ_1,
          PeriodData              => PInfo_CLK_R_EQ_1_AN_S_EQ_1,
          TestSignal              => CLK_dly,
          TestSignalName          => "CLK",
          TestDelay               => ticd_CLK,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TO_X01(( (NOT S_CLK_dly) ) OR ( (NOT R_CLK_dly) )
                            ) /= '1',
          HeaderMsg               => InstancePath & "/DFFRS",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      D_delayed := D_CLK_dly;
      CLK_delayed := CLK_dly;
      Violation := Tviol_D_CLK_R_EQ_1_AN_S_EQ_1_posedge or Tviol_R_CLK_S_EQ_1_posedge or Tviol_S_CLK_R_EQ_1_posedge or Pviol_CLK_R_EQ_1_AN_S_EQ_1 or Pviol_R or Pviol_S;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => dfftab,
        DataIn => (
               D_delayed, CLK_delayed, R_CLK_dly, S_CLK_dly));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (R_CLK_dly'last_event, tpd_R_Q, TRUE),
                 1 => (S_CLK_dly'last_event, tpd_S_Q, TRUE),
                 2 => (CLK_dly'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;

configuration CFG_DFFRS_VITAL of DFFRS is 
        for VITAL_VF
        end for; 
end CFG_DFFRS_VITAL;
----- VITAL model for cell DFFRSH -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;
LIBRARY VF1 ;
use VF1.VLOGTOVITAL_TABLES.all;

-- entity declaration --
entity DFFRSH is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_R_Q                        :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tpd_S_Q                        :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tsetup_D_CLK_noedge_posedge    :	VitalDelayType := 2.200 ns;
      thold_D_CLK_noedge_posedge     :	VitalDelayType := 2.200 ns;
      tpw_CLK_posedge 		     :	VitalDelayType := 4.400 ns;
      tpw_R_posedge 		     :	VitalDelayType := 4.400 ns;
      tpw_S_posedge 		     :	VitalDelayType := 4.400 ns;
      tperiod_CLK_posedge   	     :	VitalDelayType := 8.800 ns;
      trecovery_R_CLK_negedge_posedge :	VitalDelayType := 2.200 ns;
      thold_R_CLK_negedge_posedge     :	VitalDelayType := 2.200 ns;
      trecovery_S_CLK_negedge_posedge :	VitalDelayType := 2.200 ns;
      thold_S_CLK_negedge_posedge     :	VitalDelayType := 2.200 ns;
      ticd_CLK                        :	VitalDelayType := 0.000 ns;
      tisd_D_CLK                      :	VitalDelayType := 0.000 ns;
      tisd_R_CLK                      :	VitalDelayType := 0.000 ns;
      tisd_S_CLK                      :	VitalDelayType := 0.000 ns;
      tipd_D                          :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_R                          :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                          :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      R                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFFRSH : entity is TRUE;
end DFFRSH;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library VF1;
architecture VITAL_VF of DFFRSH is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL R_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL D_CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL R_CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL S_CLK_dly	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (R_ipd, R, tipd_R);
   VitalWireDelay (S_ipd, S, tipd_S);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   VitalSignalDelay (CLK_dly, CLK_ipd, ticd_CLK);
   VitalSignalDelay (D_CLK_dly, D_ipd, tisd_D_CLK);
   VitalSignalDelay (R_CLK_dly, R_ipd, tisd_R_CLK);
   VitalSignalDelay (S_CLK_dly, S_ipd, tisd_S_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (CLK_dly, D_CLK_dly, R_CLK_dly, S_CLK_dly)

   -- timing check results
   VARIABLE Tviol_D_CLK_R_EQ_0_AN_S_EQ_0_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_R_EQ_0_AN_S_EQ_0_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_R_CLK_S_EQ_0_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_R_CLK_S_EQ_0_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S_CLK_R_EQ_0_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S_CLK_R_EQ_0_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK_R_EQ_0_AN_S_EQ_0	: STD_ULOGIC := '0';
   VARIABLE Pviol_R			: STD_ULOGIC := '0';
   VARIABLE Pviol_S			: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK_R_EQ_0_AN_S_EQ_0	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE PInfo_R			: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE PInfo_S			: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(1 to 4);
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE R_inverted: STD_ULOGIC := 'X';
   VARIABLE S_inverted : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_R_EQ_0_AN_S_EQ_0_posedge,
          TimingData              => Tmkr_D_CLK_R_EQ_0_AN_S_EQ_0_posedge,
          TestSignal              => D_CLK_dly,
          TestSignalName          => "D",
          TestDelay               => tisd_D_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          SetupHigh               => tsetup_D_CLK_noedge_posedge,
          SetupLow                => tsetup_D_CLK_noedge_posedge,
          HoldHigh                => thold_D_CLK_noedge_posedge,
          HoldLow                 => thold_D_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(((NOT S_CLK_dly)) AND ((NOT R_CLK_dly))) /=
                            '0',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFFRSH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_R_CLK_S_EQ_0_posedge,
          TimingData              => Tmkr_R_CLK_S_EQ_0_posedge,
          TestSignal              => R_CLK_dly,
          TestSignalName          => "R",
          TestDelay               => tisd_R_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          Recovery                => trecovery_R_CLK_negedge_posedge,
          Removal                 => thold_R_CLK_negedge_posedge,
          ActiveLow               => FALSE,
          CheckEnabled            => 
                           TO_X01((NOT S_CLK_dly)) /= '0',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFFRSH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_S_CLK_R_EQ_0_posedge,
          TimingData              => Tmkr_S_CLK_R_EQ_0_posedge,
          TestSignal              => S_CLK_dly,
          TestSignalName          => "S",
          TestDelay               => tisd_S_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          Recovery                => trecovery_S_CLK_negedge_posedge,
          Removal                 => thold_S_CLK_negedge_posedge,
          ActiveLow               => FALSE,
          CheckEnabled            => 
                           TO_X01((NOT R_CLK_dly)) /= '0',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFFRSH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_S,
          PeriodData              => PInfo_S,
          TestSignal              => R_CLK_dly,
          TestSignalName          => "R",
          TestDelay               => tisd_S_CLK,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_S_posedge,
          CheckEnabled            => TRUE, 
          HeaderMsg               => InstancePath & "/DFFRSH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_R,
          PeriodData              => PInfo_R,
          TestSignal              => R_CLK_dly,
          TestSignalName          => "R",
          TestDelay               => tisd_R_CLK,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_R_posedge,
          CheckEnabled            => TRUE, 
          HeaderMsg               => InstancePath & "/DFFRSH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK_R_EQ_0_AN_S_EQ_0,
          PeriodData              => PInfo_CLK_R_EQ_0_AN_S_EQ_0,
          TestSignal              => CLK_dly,
          TestSignalName          => "CLK",
          TestDelay               => ticd_CLK,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TO_X01(( S_CLK_dly ) OR ( R_CLK_dly ) ) /= '1',
          HeaderMsg               => InstancePath & "/DFFRSH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      D_delayed := D_CLK_dly;
      CLK_delayed := CLK_dly;
      R_inverted := NOT R_CLK_dly;
      S_inverted := NOT S_CLK_dly;
      Violation := Tviol_D_CLK_R_EQ_0_AN_S_EQ_0_posedge or Tviol_R_CLK_S_EQ_0_posedge or Tviol_S_CLK_R_EQ_0_posedge or Pviol_CLK_R_EQ_0_AN_S_EQ_0 or Pviol_R or Pviol_S;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => dfftab,
        DataIn => (
               D_delayed, CLK_delayed, R_inverted, S_inverted));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (R_CLK_dly'last_event, tpd_R_Q, TRUE),
                 1 => (S_CLK_dly'last_event, tpd_S_Q, TRUE),
                 2 => (CLK_dly'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;

configuration CFG_DFFRSH_VITAL of DFFRSH is 
        for VITAL_VF
        end for; 
end CFG_DFFRSH_VITAL;
----- VITAL model for cell DFFRSS -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;

LIBRARY VF1 ;
use VF1.VLOGTOVITAL_TABLES.all;



-- entity declaration --
entity DFFRSS is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_R_Q                        :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tpd_S_Q                        :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tsetup_D_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      thold_D_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      tpw_CLK_posedge :	VitalDelayType := 4.400 ns;
      tperiod_CLK_posedge  :	VitalDelayType := 8.800 ns;
      trecovery_R_CLK_posedge_posedge :	VitalDelayType := 2.200 ns;
      thold_R_CLK_posedge_posedge :	VitalDelayType := 2.200 ns;
      trecovery_S_CLK_posedge_posedge :	VitalDelayType := 2.200 ns;
      thold_S_CLK_posedge_posedge :	VitalDelayType := 2.200 ns;
      ticd_CLK                       :	VitalDelayType := 0.000 ns;
      tisd_D_CLK                     :	VitalDelayType := 0.000 ns;
      tisd_R_CLK                     :	VitalDelayType := 0.000 ns;
      tisd_S_CLK                     :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_R                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      R                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFFRSS : entity is TRUE;
end DFFRSS;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library VF1;
architecture VITAL_VF of DFFRSS is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL R_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL D_CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL R_CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL S_CLK_dly	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (R_ipd, R, tipd_R);
   VitalWireDelay (S_ipd, S, tipd_S);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   VitalSignalDelay (CLK_dly, CLK_ipd, ticd_CLK);
   VitalSignalDelay (D_CLK_dly, D_ipd, tisd_D_CLK);
   VitalSignalDelay (R_CLK_dly, R_ipd, tisd_R_CLK);
   VitalSignalDelay (S_CLK_dly, S_ipd, tisd_S_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (CLK_dly, D_CLK_dly, R_CLK_dly, S_CLK_dly)

   -- timing check results
   VARIABLE Tviol_D_CLK_R_EQ_1_ANB_S_EQ_1_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_R_EQ_1_ANB_S_EQ_1_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_R_CLK_S_EQ_1_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_R_CLK_S_EQ_1_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S_CLK_R_EQ_1_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S_CLK_R_EQ_1_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK_R_EQ_1_ANB_S_EQ_1	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK_R_EQ_1_ANB_S_EQ_1	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 3);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);
   VARIABLE NOT_S_zd : STD_ULOGIC := '0';
   VARIABLE D_in_zd : STD_ULOGIC := '0';

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_R_EQ_1_ANB_S_EQ_1_posedge,
          TimingData              => Tmkr_D_CLK_R_EQ_1_ANB_S_EQ_1_posedge,
          TestSignal              => D_CLK_dly,
          TestSignalName          => "D",
          TestDelay               => tisd_D_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          SetupHigh               => tsetup_D_CLK_noedge_posedge,
          SetupLow                => tsetup_D_CLK_noedge_posedge,
          HoldHigh                => thold_D_CLK_noedge_posedge,
          HoldLow                 => thold_D_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((S_CLK_dly) AND (R_CLK_dly)) = '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFFRSS",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_R_CLK_S_EQ_1_posedge,
          TimingData              => Tmkr_R_CLK_S_EQ_1_posedge,
          TestSignal              => R_CLK_dly,
          TestSignalName          => "R",
          TestDelay               => tisd_R_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          Recovery                => trecovery_R_CLK_posedge_posedge,
          Removal                 => thold_R_CLK_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TO_X01(S_CLK_dly) = '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFFRSS",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_S_CLK_R_EQ_1_posedge,
          TimingData              => Tmkr_S_CLK_R_EQ_1_posedge,
          TestSignal              => S_CLK_dly,
          TestSignalName          => "S",
          TestDelay               => tisd_S_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          Recovery                => trecovery_S_CLK_posedge_posedge,
          Removal                 => thold_S_CLK_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TO_X01(R_CLK_dly) = '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFFRSS",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK_R_EQ_1_ANB_S_EQ_1,
          PeriodData              => PInfo_CLK_R_EQ_1_ANB_S_EQ_1,
          TestSignal              => CLK_dly,
          TestSignalName          => "CLK",
          TestDelay               => ticd_CLK,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TO_X01(( (S_CLK_dly) ) AND ( (R_CLK_dly) )) = '1',
          HeaderMsg               => InstancePath & "/DFFRSS",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------

        NOT_S_zd := VitalINV (S_CLK_dly);
        D_in_zd := VitalOR2 (NOT_S_zd , D_CLK_dly);

      Violation := Tviol_D_CLK_R_EQ_1_ANB_S_EQ_1_posedge or Tviol_R_CLK_S_EQ_1_posedge or Tviol_S_CLK_R_EQ_1_posedge or Pviol_CLK_R_EQ_1_ANB_S_EQ_1;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => dfftab,
        DataIn => (
               D_in_zd, CLK_dly, R_CLK_dly, '1'));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (R_CLK_dly'last_event, tpd_R_Q, TRUE),
                 1 => (S_CLK_dly'last_event, tpd_S_Q, TRUE),
                 2 => (CLK_dly'last_event, tpd_CLK_Q, TRUE)),
       Mode => VitalInertial,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;

configuration CFG_DFFRSS_VITAL of DFFRSS is 
        for VITAL_VF
        end for; 
end CFG_DFFRSS_VITAL;
----- VITAL model for cell DFFRSSH -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;

LIBRARY VF1 ;
use VF1.VLOGTOVITAL_TABLES.all;



-- entity declaration --
entity DFFRSSH is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_R_Q                        :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tpd_S_Q                        :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tsetup_D_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      thold_D_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      tpw_CLK_posedge :	VitalDelayType := 4.400 ns;
      tpw_R_posedge :	VitalDelayType := 4.400 ns;
      tperiod_CLK_posedge  :	VitalDelayType := 8.800 ns;
      trecovery_R_CLK_negedge_posedge :	VitalDelayType := 2.200 ns;
      thold_R_CLK_negedge_posedge :	VitalDelayType := 2.200 ns;
      tsetup_S_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      thold_S_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      ticd_CLK                       :	VitalDelayType := 0.000 ns;
      tisd_D_CLK                     :	VitalDelayType := 0.000 ns;
      tisd_R_CLK                     :	VitalDelayType := 0.000 ns;
      tisd_S_CLK                     :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_R                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      R                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFFRSSH : entity is TRUE;
end DFFRSSH;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library VF1;
architecture VITAL_VF of DFFRSSH is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL R_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL D_CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL R_CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL S_CLK_dly	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (R_ipd, R, tipd_R);
   VitalWireDelay (S_ipd, S, tipd_S);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   VitalSignalDelay (CLK_dly, CLK_ipd, ticd_CLK);
   VitalSignalDelay (D_CLK_dly, D_ipd, tisd_D_CLK);
   VitalSignalDelay (R_CLK_dly, R_ipd, tisd_R_CLK);
   VitalSignalDelay (S_CLK_dly, S_ipd, tisd_S_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (CLK_dly, D_CLK_dly, R_CLK_dly, S_CLK_dly)

   -- timing check results
   VARIABLE Tviol_D_CLK_R_EQ_0_ANB_S_EQ_0_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_R_EQ_0_ANB_S_EQ_0_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_R_CLK_S_EQ_0_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_R_CLK_S_EQ_0_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S_CLK_R_EQ_0_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S_CLK_R_EQ_0_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK_R_EQ_0_ANB_S_EQ_0	: STD_ULOGIC := '0';
   VARIABLE Pviol_R	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK_R_EQ_0_ANB_S_EQ_0	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE PInfo_R	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 3);
   VARIABLE R_inverted : STD_ULOGIC := 'X';
   VARIABLE S_inverted : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);
   VARIABLE D_in_zd : STD_ULOGIC := '0';


   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_R_EQ_0_ANB_S_EQ_0_posedge,
          TimingData              => Tmkr_D_CLK_R_EQ_0_ANB_S_EQ_0_posedge,
          TestSignal              => D_CLK_dly,
          TestSignalName          => "D",
          TestDelay               => tisd_D_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          SetupHigh               => tsetup_D_CLK_noedge_posedge,
          SetupLow                => tsetup_D_CLK_noedge_posedge,
          HoldHigh                => thold_D_CLK_noedge_posedge,
          HoldLow                 => thold_D_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(((NOT S_CLK_dly)) AND ((NOT R_CLK_dly))) = '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFFRSSH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_R_CLK_S_EQ_0_posedge,
          TimingData              => Tmkr_R_CLK_S_EQ_0_posedge,
          TestSignal              => R_CLK_dly,
          TestSignalName          => "R",
          TestDelay               => tisd_R_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          Recovery                => trecovery_R_CLK_negedge_posedge,
          Removal                 => thold_R_CLK_negedge_posedge,
          ActiveLow               => FALSE,
          CheckEnabled            => 
                           TO_X01((NOT S_CLK_dly)) = '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFFRSSH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_S_CLK_R_EQ_0_posedge,
          TimingData              => Tmkr_S_CLK_R_EQ_0_posedge,
          TestSignal              => S_CLK_dly,
          TestSignalName          => "S",
          TestDelay               => tisd_S_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          SetupHigh               => tsetup_S_CLK_noedge_posedge,
          SetupLow                => tsetup_S_CLK_noedge_posedge,
          HoldHigh                => thold_S_CLK_noedge_posedge,
          HoldLow                 => thold_S_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT R_CLK_dly)) = '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFFRSSH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_R,
          PeriodData              => PInfo_R,
          TestSignal              => R_CLK_dly,
          TestSignalName          => "R",
          TestDelay               => tisd_R_CLK,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_R_posedge,
          CheckEnabled            => TRUE, 
          HeaderMsg               => InstancePath & "/DFFRSSH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK_R_EQ_0_ANB_S_EQ_0,
          PeriodData              => PInfo_CLK_R_EQ_0_ANB_S_EQ_0,
          TestSignal              => CLK_dly,
          TestSignalName          => "CLK",
          TestDelay               => ticd_CLK,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TO_X01(((NOT S_CLK_dly)) AND ((NOT R_CLK_dly))) = '1',
          HeaderMsg               => InstancePath & "/DFFRSSH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------

        D_in_zd := VitalOR2 (S_CLK_dly , D_CLK_dly);

      Violation := Tviol_D_CLK_R_EQ_0_ANB_S_EQ_0_posedge or Tviol_S_CLK_R_EQ_0_posedge or Pviol_CLK_R_EQ_0_ANB_S_EQ_0 or Tviol_R_CLK_S_EQ_0_posedge or Pviol_R;
      S_inverted := (NOT S_CLK_dly);
      R_inverted := (NOT R_CLK_dly);
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => dfftab,
        DataIn => (
               D_in_zd, CLK_dly, R_inverted, '1' ));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (R_CLK_dly'last_event, tpd_R_Q, TRUE),
                 1 => (S_CLK_dly'last_event, tpd_S_Q, TRUE),
                 2 => (CLK_dly'last_event, tpd_CLK_Q, TRUE)),
       Mode => VitalInertial,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;

configuration CFG_DFFRSSH_VITAL of DFFRSSH is 
        for VITAL_VF
        end for; 
end CFG_DFFRSSH_VITAL;
----- VITAL model for cell DFFS -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;

LIBRARY VF1 ;
use VF1.VLOGTOVITAL_TABLES.all;



-- entity declaration --
entity DFFS is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_S_Q                        :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tsetup_D_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      thold_D_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      tpw_CLK_posedge         :	VitalDelayType := 4.400 ns;
      tperiod_CLK_posedge             :	VitalDelayType := 8.800 ns;
      trecovery_S_CLK_posedge_posedge :	VitalDelayType := 2.200 ns;
      thold_S_CLK_posedge_posedge    :	VitalDelayType := 2.200 ns;
      ticd_CLK                       :	VitalDelayType := 0.000 ns;
      tisd_D_CLK                     :	VitalDelayType := 0.000 ns;
      tisd_S_CLK                     :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFFS : entity is TRUE;
end DFFS;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library VF1;
architecture VITAL_VF of DFFS is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL D_CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL S_CLK_dly	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (S_ipd, S, tipd_S);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   VitalSignalDelay (CLK_dly, CLK_ipd, ticd_CLK);
   VitalSignalDelay (D_CLK_dly, D_ipd, tisd_D_CLK);
   VitalSignalDelay (S_CLK_dly, S_ipd, tisd_S_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (CLK_dly, D_CLK_dly, S_CLK_dly)

   -- timing check results
   VARIABLE Tviol_D_CLK_S_EQ_1_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_S_EQ_1_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK_S_EQ_1	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK_S_EQ_1	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 3);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_S_EQ_1_posedge,
          TimingData              => Tmkr_D_CLK_S_EQ_1_posedge,
          TestSignal              => D_CLK_dly,
          TestSignalName          => "D",
          TestDelay               => tisd_D_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          SetupHigh               => tsetup_D_CLK_noedge_posedge,
          SetupLow                => tsetup_D_CLK_noedge_posedge,
          HoldHigh                => thold_D_CLK_noedge_posedge,
          HoldLow                 => thold_D_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(S_CLK_dly) = '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFFS",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_S_CLK_posedge,
          TimingData              => Tmkr_S_CLK_posedge,
          TestSignal              => S_CLK_dly,
          TestSignalName          => "S",
          TestDelay               => tisd_S_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          Recovery                => trecovery_S_CLK_posedge_posedge,
          Removal                 => thold_S_CLK_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFFS",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK_S_EQ_1,
          PeriodData              => PInfo_CLK_S_EQ_1,
          TestSignal              => CLK_dly,
          TestSignalName          => "CLK",
          TestDelay               => ticd_CLK,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TO_X01((S_CLK_dly) ) = '1',
          HeaderMsg               => InstancePath & "/DFFS",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_S_EQ_1_posedge or Tviol_S_CLK_posedge or Pviol_CLK_S_EQ_1;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => dfftab,
        DataIn => (
               D_CLK_dly, CLK_dly, '1', S_CLK_dly));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (S_CLK_dly'last_event, tpd_S_Q, TRUE),
                 1 => (CLK_dly'last_event, tpd_CLK_Q, TRUE)),
       Mode => VitalInertial,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;

configuration CFG_DFFS_VITAL of DFFS is 
        for VITAL_VF
        end for; 
end CFG_DFFS_VITAL;
----- VITAL model for cell DFFSH -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;

LIBRARY VF1 ;
use VF1.VLOGTOVITAL_TABLES.all;



-- entity declaration --
entity DFFSH is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_S_Q                        :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tsetup_D_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      thold_D_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      tpw_CLK_posedge         :	VitalDelayType := 4.400 ns;
      tpw_S_posedge         :	VitalDelayType := 4.400 ns;
      tperiod_CLK_posedge             :	VitalDelayType := 8.800 ns;
      trecovery_S_CLK_negedge_posedge :	VitalDelayType := 2.200 ns;
      thold_S_CLK_negedge_posedge    :	VitalDelayType := 2.200 ns;
      ticd_CLK                       :	VitalDelayType := 0.000 ns;
      tisd_D_CLK                     :	VitalDelayType := 0.000 ns;
      tisd_S_CLK                     :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFFSH : entity is TRUE;
end DFFSH;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library VF1;
architecture VITAL_VF of DFFSH is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL D_CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL S_CLK_dly	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (S_ipd, S, tipd_S);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   VitalSignalDelay (CLK_dly, CLK_ipd, ticd_CLK);
   VitalSignalDelay (D_CLK_dly, D_ipd, tisd_D_CLK);
   VitalSignalDelay (S_CLK_dly, S_ipd, tisd_S_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (CLK_dly, D_CLK_dly, S_CLK_dly)

   -- timing check results
   VARIABLE Tviol_D_CLK_S_EQ_0_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_S_EQ_0_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK_S_EQ_0	: STD_ULOGIC := '0';
   VARIABLE Pviol_S	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK_S_EQ_0	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE PInfo_S	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 3);
   VARIABLE S_inverted : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_S_EQ_0_posedge,
          TimingData              => Tmkr_D_CLK_S_EQ_0_posedge,
          TestSignal              => D_CLK_dly,
          TestSignalName          => "D",
          TestDelay               => tisd_D_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          SetupHigh               => tsetup_D_CLK_noedge_posedge,
          SetupLow                => tsetup_D_CLK_noedge_posedge,
          HoldHigh                => thold_D_CLK_noedge_posedge,
          HoldLow                 => thold_D_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((S_CLK_dly)) = '0',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFFSH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_S_CLK_posedge,
          TimingData              => Tmkr_S_CLK_posedge,
          TestSignal              => S_CLK_dly,
          TestSignalName          => "S",
          TestDelay               => tisd_S_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          Recovery                => trecovery_S_CLK_negedge_posedge,
          Removal                 => thold_S_CLK_negedge_posedge,
          ActiveLow               => FALSE,
          CheckEnabled            => TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFFSH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_S,
          PeriodData              => PInfo_S,
          TestSignal              => S_CLK_dly,
          TestSignalName          => "S",
          TestDelay               => tisd_S_CLK,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_S_posedge,
          CheckEnabled            => TRUE, 
          HeaderMsg               => InstancePath & "/DFFSH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK_S_EQ_0,
          PeriodData              => PInfo_CLK_S_EQ_0,
          TestSignal              => CLK_dly,
          TestSignalName          => "CLK",
          TestDelay               => ticd_CLK,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TO_X01(S_CLK_dly ) = '0',
          HeaderMsg               => InstancePath & "/DFFSH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_S_EQ_0_posedge or Tviol_S_CLK_posedge or Pviol_CLK_S_EQ_0;
      S_inverted := (NOT S_CLK_dly);
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => dfftab,
        DataIn => (
               D_CLK_dly, CLK_dly, '1', S_inverted));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (S_CLK_dly'last_event, tpd_S_Q, TRUE),
                 1 => (CLK_dly'last_event, tpd_CLK_Q, TRUE)),
       Mode => VitalInertial,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;

configuration CFG_DFFSH_VITAL of DFFSH is 
        for VITAL_VF
        end for; 
end CFG_DFFSH_VITAL;
----- VITAL model for cell DLAT -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;

LIBRARY VF1 ;
use VF1.VLOGTOVITAL_TABLES.all;



-- entity declaration --
entity DLAT is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_D_Q                        :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tpd_LAT_Q                      :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tsetup_D_LAT_noedge_negedge    :	VitalDelayType := 2.200 ns;
      thold_D_LAT_noedge_negedge     :	VitalDelayType := 2.200 ns;
      tperiod_LAT_posedge            :	VitalDelayType := 8.800 ns;
      tpw_LAT_posedge                :	VitalDelayType := 4.400 ns;
      ticd_LAT                       :	VitalDelayType := 0.000 ns;
      tisd_D_LAT                     :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_LAT                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      LAT                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DLAT : entity is TRUE;
end DLAT;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library VF1;
architecture VITAL_VF of DLAT is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL LAT_ipd	 : STD_ULOGIC := 'X';
   SIGNAL LAT_dly	 : STD_ULOGIC := 'X';
   SIGNAL D_LAT_dly	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (LAT_ipd, LAT, tipd_LAT);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   VitalSignalDelay (LAT_dly, LAT_ipd, ticd_LAT);
   VitalSignalDelay (D_LAT_dly, D_ipd, tisd_D_LAT);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (LAT_dly, D_LAT_dly)

   -- timing check results
   VARIABLE Tviol_D_LAT_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_LAT_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_LAT	: STD_ULOGIC := '0';
   VARIABLE PInfo_LAT	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 3);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_LAT_negedge,
          TimingData              => Tmkr_D_LAT_negedge,
          TestSignal              => D_LAT_dly,
          TestSignalName          => "D",
          TestDelay               => tisd_D_LAT,
          RefSignal               => LAT_dly,
          RefSignalName          => "LAT",
          RefDelay                => ticd_LAT,
          SetupHigh               => tsetup_D_LAT_noedge_negedge,
          SetupLow                => tsetup_D_LAT_noedge_negedge,
          HoldHigh                => thold_D_LAT_noedge_negedge,
          HoldLow                 => thold_D_LAT_noedge_negedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DLAT",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_LAT,
          PeriodData              => PInfo_LAT,
          TestSignal              => LAT_dly,
          TestSignalName          => "LAT",
          TestDelay               => ticd_LAT,
          Period                  => tperiod_LAT_posedge,
          PulseWidthHigh          => tpw_LAT_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DLAT",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_LAT_negedge or Pviol_LAT;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => latchtab,
        DataIn => (
               D_LAT_dly, LAT_dly,'1','1'));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (D_LAT_dly'last_event, tpd_D_Q, TRUE),
                 1 => (LAT_dly'last_event, tpd_LAT_Q, TRUE)),
       Mode => VitalInertial,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;

configuration CFG_DLAT_VITAL of DLAT is 
        for VITAL_VF
        end for; 
end CFG_DLAT_VITAL;
----- VITAL model for cell DLATR -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;

LIBRARY VF1 ;
use VF1.VLOGTOVITAL_TABLES.all;



-- entity declaration --
entity DLATR is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_D_Q                        :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tpd_LAT_Q                      :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tpd_R_Q                        :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tsetup_D_LAT_noedge_negedge :	VitalDelayType := 2.200 ns;
      thold_D_LAT_noedge_negedge :	VitalDelayType := 2.200 ns;
      tpw_LAT_posedge         :	VitalDelayType := 4.400 ns;
      tperiod_LAT_posedge             :	VitalDelayType := 8.800 ns;
      trecovery_R_LAT_posedge_negedge :	VitalDelayType := 2.200 ns;
      thold_R_LAT_posedge_negedge    :	VitalDelayType := 2.200 ns;
      ticd_LAT                       :	VitalDelayType := 0.000 ns;
      tisd_D_LAT                     :	VitalDelayType := 0.000 ns;
      tisd_R_LAT                     :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_LAT                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_R                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      LAT                            :	in    STD_ULOGIC;
      R                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DLATR : entity is TRUE;
end DLATR;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library VF1;
architecture VITAL_VF of DLATR is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL LAT_ipd	 : STD_ULOGIC := 'X';
   SIGNAL R_ipd	 : STD_ULOGIC := 'X';
   SIGNAL LAT_dly	 : STD_ULOGIC := 'X';
   SIGNAL D_LAT_dly	 : STD_ULOGIC := 'X';
   SIGNAL R_LAT_dly	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (LAT_ipd, LAT, tipd_LAT);
   VitalWireDelay (R_ipd, R, tipd_R);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   VitalSignalDelay (LAT_dly, LAT_ipd, ticd_LAT);
   VitalSignalDelay (D_LAT_dly, D_ipd, tisd_D_LAT);
   VitalSignalDelay (R_LAT_dly, R_ipd, tisd_R_LAT);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (LAT_dly, D_LAT_dly, R_LAT_dly)

   -- timing check results
   VARIABLE Tviol_D_LAT_R_EQ_1_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_LAT_R_EQ_1_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_R_LAT_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_R_LAT_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_LAT_R_EQ_1	: STD_ULOGIC := '0';
   VARIABLE PInfo_LAT_R_EQ_1	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 3);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_LAT_R_EQ_1_negedge,
          TimingData              => Tmkr_D_LAT_R_EQ_1_negedge,
          TestSignal              => D_LAT_dly,
          TestSignalName          => "D",
          TestDelay               => tisd_D_LAT,
          RefSignal               => LAT_dly,
          RefSignalName          => "LAT",
          RefDelay                => ticd_LAT,
          SetupHigh               => tsetup_D_LAT_noedge_negedge,
          SetupLow                => tsetup_D_LAT_noedge_negedge,
          HoldHigh                => thold_D_LAT_noedge_negedge,
          HoldLow                 => thold_D_LAT_noedge_negedge,
          CheckEnabled            => 
                           TO_X01(R_LAT_dly) = '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DLATR",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_R_LAT_negedge,
          TimingData              => Tmkr_R_LAT_negedge,
          TestSignal              => R_LAT_dly,
          TestSignalName          => "R",
          TestDelay               => tisd_R_LAT,
          RefSignal               => LAT_dly,
          RefSignalName          => "LAT",
          RefDelay                => ticd_LAT,
          Recovery                => trecovery_R_LAT_posedge_negedge,
          Removal                 => thold_R_LAT_posedge_negedge,
          ActiveLow               => TRUE,
          CheckEnabled            => TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DLATR",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_LAT_R_EQ_1,
          PeriodData              => PInfo_LAT_R_EQ_1,
          TestSignal              => LAT_dly,
          TestSignalName          => "LAT",
          TestDelay               => ticd_LAT,
          Period                  => tperiod_LAT_posedge,
          PulseWidthHigh          => tpw_LAT_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TO_X01(R_LAT_dly ) = '1',
          HeaderMsg               => InstancePath & "/DLATR",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_LAT_R_EQ_1_negedge or Tviol_R_LAT_negedge or Pviol_LAT_R_EQ_1;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => latchtab,
        DataIn => (
               D_LAT_dly, LAT_dly, R_LAT_dly,'1'));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (D_LAT_dly'last_event, tpd_D_Q, TRUE),
                 1 => (LAT_dly'last_event, tpd_LAT_Q, TRUE),
                 2 => (R_LAT_dly'last_event, tpd_R_Q, TRUE)),
       Mode => VitalInertial,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;

configuration CFG_DLATR_VITAL of DLATR is 
        for VITAL_VF
        end for; 
end CFG_DLATR_VITAL;
----- VITAL model for cell DLATRH -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;

LIBRARY VF1 ;
use VF1.VLOGTOVITAL_TABLES.all;



-- entity declaration --
entity DLATRH is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_D_Q                        :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tpd_LAT_Q                      :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tpd_R_Q                        :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tsetup_D_LAT_noedge_negedge :	VitalDelayType := 2.200 ns;
      thold_D_LAT_noedge_negedge :	VitalDelayType := 2.200 ns;
      tpw_LAT_posedge         :	VitalDelayType := 4.400 ns;
      tperiod_LAT_posedge             :	VitalDelayType := 8.800 ns;
      trecovery_R_LAT_negedge_negedge :	VitalDelayType := 2.200 ns;
      thold_R_LAT_negedge_negedge    :	VitalDelayType := 2.200 ns;
      ticd_LAT                       :	VitalDelayType := 0.000 ns;
      tisd_D_LAT                     :	VitalDelayType := 0.000 ns;
      tisd_R_LAT                     :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_LAT                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_R                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      LAT                            :	in    STD_ULOGIC;
      R                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DLATRH : entity is TRUE;
end DLATRH;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library VF1;
architecture VITAL_VF of DLATRH is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL LAT_ipd	 : STD_ULOGIC := 'X';
   SIGNAL R_ipd	 : STD_ULOGIC := 'X';
   SIGNAL LAT_dly	 : STD_ULOGIC := 'X';
   SIGNAL D_LAT_dly	 : STD_ULOGIC := 'X';
   SIGNAL R_LAT_dly	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (LAT_ipd, LAT, tipd_LAT);
   VitalWireDelay (R_ipd, R, tipd_R);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   VitalSignalDelay (LAT_dly, LAT_ipd, ticd_LAT);
   VitalSignalDelay (D_LAT_dly, D_ipd, tisd_D_LAT);
   VitalSignalDelay (R_LAT_dly, R_ipd, tisd_R_LAT);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (LAT_dly, D_LAT_dly, R_LAT_dly)

   -- timing check results
   VARIABLE Tviol_D_LAT_R_EQ_0_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_LAT_R_EQ_0_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_R_LAT_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_R_LAT_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_LAT_R_EQ_0	: STD_ULOGIC := '0';
   VARIABLE PInfo_LAT_R_EQ_0	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE R_inverted : STD_ULOGIC := 'X';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 3);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_LAT_R_EQ_0_negedge,
          TimingData              => Tmkr_D_LAT_R_EQ_0_negedge,
          TestSignal              => D_LAT_dly,
          TestSignalName          => "D",
          TestDelay               => tisd_D_LAT,
          RefSignal               => LAT_dly,
          RefSignalName          => "LAT",
          RefDelay                => ticd_LAT,
          SetupHigh               => tsetup_D_LAT_noedge_negedge,
          SetupLow                => tsetup_D_LAT_noedge_negedge,
          HoldHigh                => thold_D_LAT_noedge_negedge,
          HoldLow                 => thold_D_LAT_noedge_negedge,
          CheckEnabled            => 
                           TO_X01((R_LAT_dly)) = '0',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DLATRH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_R_LAT_negedge,
          TimingData              => Tmkr_R_LAT_negedge,
          TestSignal              => R_LAT_dly,
          TestSignalName          => "R",
          TestDelay               => tisd_R_LAT,
          RefSignal               => LAT_dly,
          RefSignalName          => "LAT",
          RefDelay                => ticd_LAT,
          Recovery                => trecovery_R_LAT_negedge_negedge,
          Removal                 => thold_R_LAT_negedge_negedge,
          ActiveLow               => FALSE,
          CheckEnabled            => TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DLATRH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_LAT_R_EQ_0,
          PeriodData              => PInfo_LAT_R_EQ_0,
          TestSignal              => LAT_dly,
          TestSignalName          => "LAT",
          TestDelay               => ticd_LAT,
          Period                  => tperiod_LAT_posedge,
          PulseWidthHigh          => tpw_LAT_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TO_X01((R_LAT_dly) ) = '0',
          HeaderMsg               => InstancePath & "/DLATRH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_LAT_R_EQ_0_negedge or Tviol_R_LAT_negedge or Pviol_LAT_R_EQ_0;
      R_inverted := (NOT R_LAT_dly);
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => latchtab,
        DataIn => (
               D_LAT_dly, LAT_dly,R_inverted,'1'));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (D_LAT_dly'last_event, tpd_D_Q, TRUE),
                 1 => (LAT_dly'last_event, tpd_LAT_Q, TRUE),
                 2 => (R_LAT_dly'last_event, tpd_R_Q, TRUE)),
       Mode => VitalInertial,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;

configuration CFG_DLATRH_VITAL of DLATRH is 
        for VITAL_VF
        end for; 
end CFG_DLATRH_VITAL;
----- VITAL model for cell DLATRS -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;

LIBRARY VF1 ;
use VF1.VLOGTOVITAL_TABLES.all;



-- entity declaration --
entity DLATRS is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_D_Q                        :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tpd_LAT_Q                      :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tpd_R_Q                        :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tpd_S_Q                        :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tsetup_D_LAT_noedge_negedge :	VitalDelayType := 2.200 ns;
      thold_D_LAT_noedge_negedge :	VitalDelayType := 2.200 ns;
      tpw_LAT_posedge :	VitalDelayType := 4.400 ns;
      tpw_R_negedge :	VitalDelayType := 4.400 ns;
      tpw_S_negedge :	VitalDelayType := 4.400 ns;
      tperiod_LAT_posedge  :	VitalDelayType := 8.800 ns;
      trecovery_R_LAT_posedge_negedge :	VitalDelayType := 2.200 ns;
      thold_R_LAT_posedge_negedge :	VitalDelayType := 2.200 ns;
      trecovery_S_LAT_posedge_negedge :	VitalDelayType := 2.200 ns;
      thold_S_LAT_posedge_negedge :	VitalDelayType := 2.200 ns;
      ticd_LAT                       :	VitalDelayType := 0.000 ns;
      tisd_D_LAT                     :	VitalDelayType := 0.000 ns;
      tisd_R_LAT                     :	VitalDelayType := 0.000 ns;
      tisd_S_LAT                     :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_LAT                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_R                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      LAT                            :	in    STD_ULOGIC;
      R                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DLATRS : entity is TRUE;
end DLATRS;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library VF1;
architecture VITAL_VF of DLATRS is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL LAT_ipd	 : STD_ULOGIC := 'X';
   SIGNAL R_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S_ipd	 : STD_ULOGIC := 'X';
   SIGNAL LAT_dly	 : STD_ULOGIC := 'X';
   SIGNAL D_LAT_dly	 : STD_ULOGIC := 'X';
   SIGNAL R_LAT_dly	 : STD_ULOGIC := 'X';
   SIGNAL S_LAT_dly	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (LAT_ipd, LAT, tipd_LAT);
   VitalWireDelay (R_ipd, R, tipd_R);
   VitalWireDelay (S_ipd, S, tipd_S);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   VitalSignalDelay (LAT_dly, LAT_ipd, ticd_LAT);
   VitalSignalDelay (D_LAT_dly, D_ipd, tisd_D_LAT);
   VitalSignalDelay (R_LAT_dly, R_ipd, tisd_R_LAT);
   VitalSignalDelay (S_LAT_dly, S_ipd, tisd_S_LAT);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (LAT_dly, D_LAT_dly, R_LAT_dly, S_LAT_dly)

   -- timing check results
   VARIABLE Tviol_D_LAT_R_EQ_1_ANB_S_EQ_1_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_LAT_R_EQ_1_ANB_S_EQ_1_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_R_LAT_S_EQ_1_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_R_LAT_S_EQ_1_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S_LAT_R_EQ_1_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S_LAT_R_EQ_1_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_LAT_R_EQ_1_ANB_S_EQ_1	: STD_ULOGIC := '0';
   VARIABLE Pviol_R	: STD_ULOGIC := '0';
   VARIABLE Pviol_S	: STD_ULOGIC := '0';
   VARIABLE PInfo_LAT_R_EQ_1_ANB_S_EQ_1	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE PInfo_R	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE PInfo_S	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 3);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);
   VARIABLE D_in_zd : STD_ULOGIC := '0';
   VARIABLE NOT_S_zd : STD_ULOGIC := '0';

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_LAT_R_EQ_1_ANB_S_EQ_1_negedge,
          TimingData              => Tmkr_D_LAT_R_EQ_1_ANB_S_EQ_1_negedge,
          TestSignal              => D_LAT_dly,
          TestSignalName          => "D",
          TestDelay               => tisd_D_LAT,
          RefSignal               => LAT_dly,
          RefSignalName          => "LAT",
          RefDelay                => ticd_LAT,
          SetupHigh               => tsetup_D_LAT_noedge_negedge,
          SetupLow                => tsetup_D_LAT_noedge_negedge,
          HoldHigh                => thold_D_LAT_noedge_negedge,
          HoldLow                 => thold_D_LAT_noedge_negedge,
          CheckEnabled            => 
                           TO_X01((S_LAT_dly) AND (R_LAT_dly)) = '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DLATRS",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_R_LAT_S_EQ_1_negedge,
          TimingData              => Tmkr_R_LAT_S_EQ_1_negedge,
          TestSignal              => R_LAT_dly,
          TestSignalName          => "R",
          TestDelay               => tisd_R_LAT,
          RefSignal               => LAT_dly,
          RefSignalName          => "LAT",
          RefDelay                => ticd_LAT,
          Recovery                => trecovery_R_LAT_posedge_negedge,
          Removal                 => thold_R_LAT_posedge_negedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TO_X01(S_LAT_dly) = '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DLATRS",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_S_LAT_R_EQ_1_negedge,
          TimingData              => Tmkr_S_LAT_R_EQ_1_negedge,
          TestSignal              => S_LAT_dly,
          TestSignalName          => "S",
          TestDelay               => tisd_S_LAT,
          RefSignal               => LAT_dly,
          RefSignalName          => "LAT",
          RefDelay                => ticd_LAT,
          Recovery                => trecovery_S_LAT_posedge_negedge,
          Removal                 => thold_S_LAT_posedge_negedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TO_X01(R_LAT_dly) = '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DLATRS",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_S,
          PeriodData              => PInfo_S,
          TestSignal              => S_LAT_dly,
          TestSignalName          => "S",
          TestDelay               => tisd_S_LAT,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_S_negedge,
          CheckEnabled            => TRUE, 
          HeaderMsg               => InstancePath & "/DLATRS",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_R,
          PeriodData              => PInfo_R,
          TestSignal              => R_LAT_dly,
          TestSignalName          => "R",
          TestDelay               => tisd_R_LAT,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_R_negedge,
          CheckEnabled            => TRUE, 
          HeaderMsg               => InstancePath & "/DLATRS",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_LAT_R_EQ_1_ANB_S_EQ_1,
          PeriodData              => PInfo_LAT_R_EQ_1_ANB_S_EQ_1,
          TestSignal              => LAT_dly,
          TestSignalName          => "LAT",
          TestDelay               => ticd_LAT,
          Period                  => tperiod_LAT_posedge,
          PulseWidthHigh          => tpw_LAT_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TO_X01(( S_LAT_dly ) AND ( R_LAT_dly ) ) = '1',
          HeaderMsg               => InstancePath & "/DLATRS",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------

        NOT_S_zd := VitalINV (S_LAT_dly);
        D_in_zd := VitalOR2 (NOT_S_zd , D_LAT_dly);

      Violation := Tviol_D_LAT_R_EQ_1_ANB_S_EQ_1_negedge or Tviol_S_LAT_R_EQ_1_negedge or Pviol_LAT_R_EQ_1_ANB_S_EQ_1 or Tviol_R_LAT_S_EQ_1_negedge;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => latchtab,
        DataIn => (
               D_LAT_dly, LAT_dly, R_LAT_dly, S_LAT_dly));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (D_LAT_dly'last_event, tpd_D_Q, TRUE),
                 1 => (LAT_dly'last_event, tpd_LAT_Q, TRUE),
                 2 => (R_LAT_dly'last_event, tpd_R_Q, TRUE),
                 3 => (S_LAT_dly'last_event, tpd_S_Q, TRUE)),
       Mode => VitalInertial,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;

configuration CFG_DLATRS_VITAL of DLATRS is 
        for VITAL_VF
        end for; 
end CFG_DLATRS_VITAL;
----- VITAL model for cell DLATRSH -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;

LIBRARY VF1 ;
use VF1.VLOGTOVITAL_TABLES.all;



-- entity declaration --
entity DLATRSH is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_D_Q                        :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tpd_LAT_Q                      :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tpd_R_Q                        :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tpd_S_Q                        :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tsetup_D_LAT_noedge_negedge :	VitalDelayType := 2.200 ns;
      thold_D_LAT_noedge_negedge :	VitalDelayType := 2.200 ns;
      tpw_LAT_posedge :	VitalDelayType := 4.400 ns;
      tpw_R_posedge :	VitalDelayType := 4.400 ns;
      tpw_S_posedge :	VitalDelayType := 4.400 ns;
      tperiod_LAT_posedge  :	VitalDelayType := 8.800 ns;
      trecovery_R_LAT_negedge_negedge :	VitalDelayType := 2.200 ns;
      thold_R_LAT_negedge_negedge     :	VitalDelayType := 2.200 ns;
      trecovery_S_LAT_negedge_negedge :	VitalDelayType := 2.200 ns;
      thold_S_LAT_negedge_negedge     :	VitalDelayType := 2.200 ns;
      ticd_LAT                       :	VitalDelayType := 0.000 ns;
      tisd_D_LAT                     :	VitalDelayType := 0.000 ns;
      tisd_R_LAT                     :	VitalDelayType := 0.000 ns;
      tisd_S_LAT                     :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_LAT                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_R                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      LAT                            :	in    STD_ULOGIC;
      R                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DLATRSH : entity is TRUE;
end DLATRSH;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library VF1;
architecture VITAL_VF of DLATRSH is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL LAT_ipd	 : STD_ULOGIC := 'X';
   SIGNAL R_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S_ipd	 : STD_ULOGIC := 'X';
   SIGNAL LAT_dly	 : STD_ULOGIC := 'X';
   SIGNAL D_LAT_dly	 : STD_ULOGIC := 'X';
   SIGNAL R_LAT_dly	 : STD_ULOGIC := 'X';
   SIGNAL S_LAT_dly	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (LAT_ipd, LAT, tipd_LAT);
   VitalWireDelay (R_ipd, R, tipd_R);
   VitalWireDelay (S_ipd, S, tipd_S);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   VitalSignalDelay (LAT_dly, LAT_ipd, ticd_LAT);
   VitalSignalDelay (D_LAT_dly, D_ipd, tisd_D_LAT);
   VitalSignalDelay (R_LAT_dly, R_ipd, tisd_R_LAT);
   VitalSignalDelay (S_LAT_dly, S_ipd, tisd_S_LAT);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (LAT_dly, D_LAT_dly, R_LAT_dly, S_LAT_dly)

   -- timing check results
   VARIABLE Tviol_D_LAT_R_EQ_0_ANB_S_EQ_0_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_LAT_R_EQ_0_ANB_S_EQ_0_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_R_LAT_S_EQ_0_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_R_LAT_S_EQ_0_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S_LAT_R_EQ_0_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S_LAT_R_EQ_0_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_LAT_R_EQ_0_ANB_S_EQ_0	: STD_ULOGIC := '0';
   VARIABLE Pviol_R : STD_ULOGIC := '0';
   VARIABLE Pviol_S : STD_ULOGIC := '0';
   VARIABLE PInfo_LAT_R_EQ_0_ANB_S_EQ_0	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE PInfo_R	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE PInfo_S	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 3);
   VARIABLE R_inverted : STD_ULOGIC := 'X';
   VARIABLE S_inverted : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);
   VARIABLE D_in_zd : STD_ULOGIC := '0';

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_LAT_R_EQ_0_ANB_S_EQ_0_negedge,
          TimingData              => Tmkr_D_LAT_R_EQ_0_ANB_S_EQ_0_negedge,
          TestSignal              => D_LAT_dly,
          TestSignalName          => "D",
          TestDelay               => tisd_D_LAT,
          RefSignal               => LAT_dly,
          RefSignalName          => "LAT",
          RefDelay                => ticd_LAT,
          SetupHigh               => tsetup_D_LAT_noedge_negedge,
          SetupLow                => tsetup_D_LAT_noedge_negedge,
          HoldHigh                => thold_D_LAT_noedge_negedge,
          HoldLow                 => thold_D_LAT_noedge_negedge,
          CheckEnabled            => 
                           TO_X01(((NOT S_LAT_dly)) AND ((NOT R_LAT_dly))) = '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DLATRSH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_R_LAT_S_EQ_0_negedge,
          TimingData              => Tmkr_R_LAT_S_EQ_0_negedge,
          TestSignal              => R_LAT_dly,
          TestSignalName          => "R",
          TestDelay               => tisd_R_LAT,
          RefSignal               => LAT_dly,
          RefSignalName          => "LAT",
          RefDelay                => ticd_LAT,
          Recovery                => trecovery_R_LAT_negedge_negedge,
          Removal                 => thold_R_LAT_negedge_negedge,
          ActiveLow               => FALSE,
          CheckEnabled            => 
                           TO_X01(S_LAT_dly) = '0',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DLATRSH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_S_LAT_R_EQ_0_negedge,
          TimingData              => Tmkr_S_LAT_R_EQ_0_negedge,
          TestSignal              => S_LAT_dly,
          TestSignalName          => "S",
          TestDelay               => tisd_S_LAT,
          RefSignal               => LAT_dly,
          RefSignalName          => "LAT",
          RefDelay                => ticd_LAT,
          Recovery                => trecovery_S_LAT_negedge_negedge,
          Removal                 => thold_S_LAT_negedge_negedge,
          ActiveLow               => FALSE,
          CheckEnabled            => 
                           TO_X01(R_LAT_dly) = '0',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DLATRSH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_S,
          PeriodData              => PInfo_S,
          TestSignal              => S_LAT_dly,
          TestSignalName          => "S",
          TestDelay               => tisd_S_LAT,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_S_posedge,
          CheckEnabled            => TRUE, 
          HeaderMsg               => InstancePath & "/DLATRSH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_R,
          PeriodData              => PInfo_R,
          TestSignal              => R_LAT_dly,
          TestSignalName          => "R",
          TestDelay               => tisd_R_LAT,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_R_posedge,
          CheckEnabled            => TRUE, 
          HeaderMsg               => InstancePath & "/DLATRSH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_LAT_R_EQ_0_ANB_S_EQ_0,
          PeriodData              => PInfo_LAT_R_EQ_0_ANB_S_EQ_0,
          TestSignal              => LAT_dly,
          TestSignalName          => "LAT",
          TestDelay               => ticd_LAT,
          Period                  => tperiod_LAT_posedge,
          PulseWidthHigh          => tpw_LAT_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TO_X01(((NOT S_LAT_dly)) AND ((NOT R_LAT_dly))) = '1',
          HeaderMsg               => InstancePath & "/DLATRSH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------

        D_in_zd := VitalOR2 (S_LAT_dly , D_LAT_dly);

      Violation := Tviol_D_LAT_R_EQ_0_ANB_S_EQ_0_negedge or Tviol_R_LAT_S_EQ_0_negedge or Tviol_S_LAT_R_EQ_0_negedge or Pviol_LAT_R_EQ_0_ANB_S_EQ_0 or Pviol_R or Pviol_S;
      S_inverted := (NOT S_LAT_dly);
      R_inverted := (NOT R_LAT_dly);
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => latchtab,
        DataIn => (
               D_LAT_dly, LAT_dly, R_inverted, S_inverted));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (D_LAT_dly'last_event, tpd_D_Q, TRUE),
                 1 => (LAT_dly'last_event, tpd_LAT_Q, TRUE),
                 2 => (R_LAT_dly'last_event, tpd_R_Q, TRUE),
                 3 => (S_LAT_dly'last_event, tpd_S_Q, TRUE)),
       Mode => VitalInertial,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;

configuration CFG_DLATRSH_VITAL of DLATRSH is 
        for VITAL_VF
        end for; 
end CFG_DLATRSH_VITAL;
----- VITAL model for cell DLATS -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;

LIBRARY VF1 ;
use VF1.VLOGTOVITAL_TABLES.all;



-- entity declaration --
entity DLATS is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_D_Q                        :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tpd_LAT_Q                      :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tpd_S_Q                        :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tsetup_D_LAT_noedge_negedge :	VitalDelayType := 2.200 ns;
      thold_D_LAT_noedge_negedge :	VitalDelayType := 2.200 ns;
      tpw_LAT_posedge         :	VitalDelayType := 4.400 ns;
      tperiod_LAT_posedge             :	VitalDelayType := 8.800 ns;
      trecovery_S_LAT_posedge_negedge :	VitalDelayType := 2.200 ns;
      thold_S_LAT_posedge_negedge    :	VitalDelayType := 2.200 ns;
      ticd_LAT                       :	VitalDelayType := 0.000 ns;
      tisd_D_LAT                     :	VitalDelayType := 0.000 ns;
      tisd_S_LAT                     :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_LAT                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      LAT                            :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DLATS : entity is TRUE;
end DLATS;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library VF1;
architecture VITAL_VF of DLATS is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL LAT_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S_ipd	 : STD_ULOGIC := 'X';
   SIGNAL LAT_dly	 : STD_ULOGIC := 'X';
   SIGNAL D_LAT_dly	 : STD_ULOGIC := 'X';
   SIGNAL S_LAT_dly	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (LAT_ipd, LAT, tipd_LAT);
   VitalWireDelay (S_ipd, S, tipd_S);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   VitalSignalDelay (LAT_dly, LAT_ipd, ticd_LAT);
   VitalSignalDelay (D_LAT_dly, D_ipd, tisd_D_LAT);
   VitalSignalDelay (S_LAT_dly, S_ipd, tisd_S_LAT);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (LAT_dly, D_LAT_dly, S_LAT_dly)

   -- timing check results
   VARIABLE Tviol_D_LAT_S_EQ_1_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_LAT_S_EQ_1_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S_LAT_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S_LAT_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_LAT_S_EQ_1	: STD_ULOGIC := '0';
   VARIABLE PInfo_LAT_S_EQ_1	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 3);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_LAT_S_EQ_1_negedge,
          TimingData              => Tmkr_D_LAT_S_EQ_1_negedge,
          TestSignal              => D_LAT_dly,
          TestSignalName          => "D",
          TestDelay               => tisd_D_LAT,
          RefSignal               => LAT_dly,
          RefSignalName          => "LAT",
          RefDelay                => ticd_LAT,
          SetupHigh               => tsetup_D_LAT_noedge_negedge,
          SetupLow                => tsetup_D_LAT_noedge_negedge,
          HoldHigh                => thold_D_LAT_noedge_negedge,
          HoldLow                 => thold_D_LAT_noedge_negedge,
          CheckEnabled            => 
                           TO_X01(S_LAT_dly) = '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DLATS",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_S_LAT_negedge,
          TimingData              => Tmkr_S_LAT_negedge,
          TestSignal              => S_LAT_dly,
          TestSignalName          => "S",
          TestDelay               => tisd_S_LAT,
          RefSignal               => LAT_dly,
          RefSignalName          => "LAT",
          RefDelay                => ticd_LAT,
          Recovery                => trecovery_S_LAT_posedge_negedge,
          Removal                 => thold_S_LAT_posedge_negedge,
          ActiveLow               => TRUE,
          CheckEnabled            => TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DLATS",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_LAT_S_EQ_1,
          PeriodData              => PInfo_LAT_S_EQ_1,
          TestSignal              => LAT_dly,
          TestSignalName          => "LAT",
          TestDelay               => ticd_LAT,
          Period                  => tperiod_LAT_posedge,
          PulseWidthHigh          => tpw_LAT_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TO_X01(S_LAT_dly ) = '1',
          HeaderMsg               => InstancePath & "/DLATS",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_LAT_S_EQ_1_negedge or Tviol_S_LAT_negedge or Pviol_LAT_S_EQ_1;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => latchtab,
        DataIn => (
               D_LAT_dly, LAT_dly,'1', S_LAT_dly));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (D_LAT_dly'last_event, tpd_D_Q, TRUE),
                 1 => (LAT_dly'last_event, tpd_LAT_Q, TRUE),
                 2 => (S_LAT_dly'last_event, tpd_S_Q, TRUE)),
       Mode => VitalInertial,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;

configuration CFG_DLATS_VITAL of DLATS is 
        for VITAL_VF
        end for; 
end CFG_DLATS_VITAL;
----- VITAL model for cell DLATSH -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;

LIBRARY VF1 ;
use VF1.VLOGTOVITAL_TABLES.all;



-- entity declaration --
entity DLATSH is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_D_Q                        :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tpd_LAT_Q                      :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tpd_S_Q                        :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tsetup_D_LAT_noedge_negedge :	VitalDelayType := 2.200 ns;
      thold_D_LAT_noedge_negedge :	VitalDelayType := 2.200 ns;
      tpw_LAT_posedge         :	VitalDelayType := 4.400 ns;
      tpw_S_posedge         :	VitalDelayType := 4.400 ns;
      tperiod_LAT_posedge             :	VitalDelayType := 8.800 ns;
      trecovery_S_LAT_negedge_negedge :	VitalDelayType := 2.200 ns;
      thold_S_LAT_negedge_negedge    :	VitalDelayType := 2.200 ns;
      ticd_LAT                       :	VitalDelayType := 0.000 ns;
      tisd_D_LAT                     :	VitalDelayType := 0.000 ns;
      tisd_S_LAT                     :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_LAT                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      LAT                            :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DLATSH : entity is TRUE;
end DLATSH;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library VF1;
architecture VITAL_VF of DLATSH is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL LAT_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S_ipd	 : STD_ULOGIC := 'X';
   SIGNAL LAT_dly	 : STD_ULOGIC := 'X';
   SIGNAL D_LAT_dly	 : STD_ULOGIC := 'X';
   SIGNAL S_LAT_dly	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (LAT_ipd, LAT, tipd_LAT);
   VitalWireDelay (S_ipd, S, tipd_S);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   VitalSignalDelay (LAT_dly, LAT_ipd, ticd_LAT);
   VitalSignalDelay (D_LAT_dly, D_ipd, tisd_D_LAT);
   VitalSignalDelay (S_LAT_dly, S_ipd, tisd_S_LAT);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (LAT_dly, D_LAT_dly, S_LAT_dly)

   -- timing check results
   VARIABLE Tviol_D_LAT_S_EQ_0_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_LAT_S_EQ_0_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S_LAT_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S_LAT_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_LAT_S_EQ_0	: STD_ULOGIC := '0';
   VARIABLE Pviol_S	: STD_ULOGIC := '0';
   VARIABLE PInfo_LAT_S_EQ_0	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE PInfo_S	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 3);
   VARIABLE S_inverted : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_LAT_S_EQ_0_negedge,
          TimingData              => Tmkr_D_LAT_S_EQ_0_negedge,
          TestSignal              => D_LAT_dly,
          TestSignalName          => "D",
          TestDelay               => tisd_D_LAT,
          RefSignal               => LAT_dly,
          RefSignalName          => "LAT",
          RefDelay                => ticd_LAT,
          SetupHigh               => tsetup_D_LAT_noedge_negedge,
          SetupLow                => tsetup_D_LAT_noedge_negedge,
          HoldHigh                => thold_D_LAT_noedge_negedge,
          HoldLow                 => thold_D_LAT_noedge_negedge,
          CheckEnabled            => 
                           TO_X01((S_LAT_dly)) = '0',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DLATSH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_S_LAT_negedge,
          TimingData              => Tmkr_S_LAT_negedge,
          TestSignal              => S_LAT_dly,
          TestSignalName          => "S",
          TestDelay               => tisd_S_LAT,
          RefSignal               => LAT_dly,
          RefSignalName          => "LAT",
          RefDelay                => ticd_LAT,
          Recovery                => trecovery_S_LAT_negedge_negedge,
          Removal                 => thold_S_LAT_negedge_negedge,
          ActiveLow               => FALSE,
          CheckEnabled            => TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DLATSH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_S,
          PeriodData              => PInfo_S,
          TestSignal              => S_LAT_dly,
          TestSignalName          => "S",
          TestDelay               => tisd_S_LAT,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_S_posedge,
          CheckEnabled            => TRUE, 
          HeaderMsg               => InstancePath & "/DLATSH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_LAT_S_EQ_0,
          PeriodData              => PInfo_LAT_S_EQ_0,
          TestSignal              => LAT_dly,
          TestSignalName          => "LAT",
          TestDelay               => ticd_LAT,
          Period                  => tperiod_LAT_posedge,
          PulseWidthHigh          => tpw_LAT_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TO_X01((S_LAT_dly) ) = '0',
          HeaderMsg               => InstancePath & "/DLATSH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_LAT_S_EQ_0_negedge or Tviol_S_LAT_negedge or Pviol_LAT_S_EQ_0 or Pviol_S;
      S_inverted := (NOT S_LAT_dly);
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => latchtab,
        DataIn => (
               D_LAT_dly, LAT_dly, '1',S_inverted));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (D_LAT_dly'last_event, tpd_D_Q, TRUE),
                 1 => (LAT_dly'last_event, tpd_LAT_Q, TRUE),
                 2 => (S_LAT_dly'last_event, tpd_S_Q, TRUE)),
       Mode => VitalInertial,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;

configuration CFG_DLATSH_VITAL of DLATSH is 
        for VITAL_VF
        end for; 
end CFG_DLATSH_VITAL;
----- VITAL model for cell ENOR -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity ENOR is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_I0_O                       :	VitalDelayType01 := (1.250 ns, 1.250 ns);
      tpd_I1_O                       :	VitalDelayType01 := (1.250 ns, 1.250 ns);
      tipd_I0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      I0                             :	in    STD_ULOGIC;
      I1                             :	in    STD_ULOGIC;
      O                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of ENOR : entity is TRUE;
end ENOR;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library VF1;
--use VF1.VTABLES.all;
architecture VITAL_VF of ENOR is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL I0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I1_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (I0_ipd, I0, tipd_I0);
   VitalWireDelay (I1_ipd, I1, tipd_I1);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (I0_ipd, I1_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS O_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE O_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      O_zd := ((NOT I1_ipd)) AND ((NOT I0_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => O,
       GlitchData => O_GlitchData,
       OutSignalName => "O",
       OutTemp => O_zd,
       Paths => (0 => (I0_ipd'last_event, tpd_I0_O, TRUE),
                 1 => (I1_ipd'last_event, tpd_I1_O, TRUE)),
       Mode => VitalInertial,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;

configuration CFG_ENOR_VITAL of ENOR is 
        for VITAL_VF
        end for; 
end CFG_ENOR_VITAL;
----- VITAL model for cell EQ22 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity EQ22 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_A0_O                       :	VitalDelayType01 := (1.800 ns, 1.800 ns);
      tpd_A1_O                       :	VitalDelayType01 := (1.800 ns, 1.800 ns);
      tpd_B0_O                       :	VitalDelayType01 := (1.800 ns, 1.800 ns);
      tpd_B1_O                       :	VitalDelayType01 := (1.800 ns, 1.800 ns);
      tipd_A0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_A1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A0                             :	in    STD_ULOGIC;
      A1                             :	in    STD_ULOGIC;
      B0                             :	in    STD_ULOGIC;
      B1                             :	in    STD_ULOGIC;
      O                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of EQ22 : entity is TRUE;
end EQ22;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_VF of EQ22 is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL A0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL A1_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B1_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A0_ipd, A0, tipd_A0);
   VitalWireDelay (A1_ipd, A1, tipd_A1);
   VitalWireDelay (B0_ipd, B0, tipd_B0);
   VitalWireDelay (B1_ipd, B1, tipd_B1);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A0_ipd, A1_ipd, B0_ipd, B1_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS O_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE O_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      O_zd :=
       ((NOT ((B1_ipd) XOR (A1_ipd)))) AND ((NOT ((B0_ipd) XOR (A0_ipd))));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => O,
       GlitchData => O_GlitchData,
       OutSignalName => "O",
       OutTemp => O_zd,
       Paths => (0 => (A0_ipd'last_event, tpd_A0_O, TRUE),
                 1 => (A1_ipd'last_event, tpd_A1_O, TRUE),
                 2 => (B0_ipd'last_event, tpd_B0_O, TRUE),
                 3 => (B1_ipd'last_event, tpd_B1_O, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;

configuration CFG_EQ22_VITAL of EQ22 is 
        for VITAL_VF
        end for; 
end CFG_EQ22_VITAL;
----- VITAL model for cell GND -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity GND is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True);

   port(
      X                              :	out   STD_ULOGIC := '0');
attribute VITAL_LEVEL0 of GND : entity is TRUE;
end GND;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library VF1;
architecture VITAL_VF of GND is
   attribute VITAL_LEVEL0 of VITAL_VF : architecture is TRUE;

	SIGNAL SUPPLY0    :   STD_ULOGIC := '0';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   --  empty
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------

Inst1 : VitalBUF (X,SUPPLY0);

end VITAL_VF;

configuration CFG_GND_VITAL of GND is 
        for VITAL_VF
        end for; 
end CFG_GND_VITAL;
----- VITAL model for cell GSRBUF -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity GSRBUF is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_SRI_O                       :	VitalDelayType01 := (1.25 ns, 1.25 ns);
      tipd_SRI                        :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      SRI                             :	in    STD_ULOGIC;
      O                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of GSRBUF : entity is TRUE;
end GSRBUF;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library VF1;
architecture VITAL_VF of GSRBUF is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL SRI_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (SRI_ipd, SRI, tipd_SRI);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (SRI_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS O_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE O_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      O_zd := TO_X01(SRI_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => O,
       GlitchData => O_GlitchData,
       OutSignalName => "O",
       OutTemp => O_zd,
       Paths => (0 => (SRI_ipd'last_event, tpd_SRI_O, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;

configuration CFG_GSRBUF_VITAL of GSRBUF is 
        for VITAL_VF
        end for; 
end CFG_GSRBUF_VITAL;
----- VITAL model for cell IBUF -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity IBUF is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_I0_O                       :	VitalDelayType01 := ( 0.64 ns, 0.64 ns);
      tipd_I0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      I0                             :	in    STD_ULOGIC;
      O                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of IBUF : entity is TRUE;
end IBUF;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library VF1;
-- -- use VF1.VTABLES.all;
architecture VITAL_VF of IBUF is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL I0_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (I0_ipd, I0, tipd_I0);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (I0_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS O_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE O_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      O_zd := TO_X01(I0_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => O,
       GlitchData => O_GlitchData,
       OutSignalName => "O",
       OutTemp => O_zd,
       Paths => (0 => (I0_ipd'last_event, tpd_I0_O, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;

configuration CFG_IBUF_VITAL of IBUF is 
        for VITAL_VF
        end for; 
end CFG_IBUF_VITAL;
----- VITAL model for cell INV -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity INV is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_I0_O                       :	VitalDelayType01 := (1.25 ns, 1.25 ns);
      tipd_I0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      I0                             :	in    STD_ULOGIC;
      O                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of INV : entity is TRUE;
end INV;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library VF1;
architecture VITAL_VF of INV is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL I0_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (I0_ipd, I0, tipd_I0);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (I0_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS O_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE O_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      O_zd := (NOT I0_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => O,
       GlitchData => O_GlitchData,
       OutSignalName => "O",
       OutTemp => O_zd,
       Paths => (0 => (I0_ipd'last_event, tpd_I0_O, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;

configuration CFG_INV_VITAL of INV is 
        for VITAL_VF
        end for; 
end CFG_INV_VITAL;
----- VITAL model for cell INVTH -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;
library VF1;
use VF1.all;


-- entity declaration --
entity INVTH is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_OE_O                       :	VitalDelayType01z := 
               (0.640 ns, 0.640 ns, 0.640 ns, 0.640 ns, 0.640 ns, 0.640 ns);
      tpd_I0_O                       :	VitalDelayType01 := (0.640 ns, 0.640 ns);
      tipd_I0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_OE                        :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      I0                             :	in    STD_ULOGIC;
      OE                             :	in    STD_ULOGIC;
      O                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of INVTH : entity is TRUE;
end INVTH;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library VF1;
architecture VITAL_VF of INVTH is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL I0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL OE_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (I0_ipd, I0, tipd_I0);
   VitalWireDelay (OE_ipd, OE, tipd_OE);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (I0_ipd, OE_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS O_zd : STD_LOGIC is Results(1);
   -- output glitch detection variables
   VARIABLE O_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      O_zd := VitalBUFIF0 (data => (NOT I0_ipd),
              enable => (NOT OE_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01Z (
       OutSignal => O,
       GlitchData => O_GlitchData,
       OutSignalName => "O",
       OutTemp => O_zd,
       Paths => (0 => (OE_ipd'last_event, VitalExtendToFillDelay(tpd_OE_O), TRUE),
                 1 => (I0_ipd'last_event, VitalExtendToFillDelay(tpd_I0_O), TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING,
       OutputMap => "UX01ZWLH-");

end process;
end VITAL_VF;

configuration CFG_INVTH_VITAL of INVTH is 
        for VITAL_VF
        end for; 
end CFG_INVTH_VITAL;
----- VITAL model for cell INVTL -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;
library VF1;
use VF1.all;


-- entity declaration --
entity INVTL is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_OE_O                       :	VitalDelayType01z := 
               (0.640 ns, 0.640 ns, 0.640 ns, 0.640 ns, 0.640 ns, 0.640 ns);
      tpd_I0_O                       :	VitalDelayType01 := (0.640 ns, 0.640 ns);
      tipd_I0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_OE                        :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      I0                             :	in    STD_ULOGIC;
      OE                             :	in    STD_ULOGIC;
      O                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of INVTL : entity is TRUE;
end INVTL;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library VF1;
architecture VITAL_VF of INVTL is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL I0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL OE_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (I0_ipd, I0, tipd_I0);
   VitalWireDelay (OE_ipd, OE, tipd_OE);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (I0_ipd, OE_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS O_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE O_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      O_zd := VitalBUFIF0 (data => (NOT I0_ipd),
              enable => OE_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01Z (
       OutSignal => O,
       GlitchData => O_GlitchData,
       OutSignalName => "O",
       OutTemp => O_zd,
       Paths => (0 => (OE_ipd'last_event, VitalExtendToFillDelay(tpd_OE_O), TRUE),
                 1 => (I0_ipd'last_event, VitalExtendToFillDelay(tpd_I0_O), TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING,
       OutputMap => "UX01ZWLH-");

end process;
end VITAL_VF;

configuration CFG_INVTL_VITAL of INVTL is 
        for VITAL_VF
        end for; 
end CFG_INVTL_VITAL;

----- VITAL model for cell JKFF -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;

LIBRARY VF1 ;
use VF1.VLOGTOVITAL_TABLES.all;



-- entity declaration --
entity JKFF is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_CLK_Q                      :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tsetup_J_CLK_noedge_posedge    :	VitalDelayType := 2.200 ns;
      thold_J_CLK_noedge_posedge     :	VitalDelayType := 2.200 ns;
      tsetup_K_CLK_noedge_posedge    :	VitalDelayType := 2.200 ns;
      thold_K_CLK_noedge_posedge     :	VitalDelayType := 2.200 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 8.800 ns;
      tpw_CLK_posedge                :	VitalDelayType := 4.400 ns;
      ticd_CLK                       :	VitalDelayType := 0.000 ns;
      tisd_J_CLK                     :	VitalDelayType := 0.000 ns;
      tisd_K_CLK                     :	VitalDelayType := 0.000 ns;
      tipd_J                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_K                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      J                              :	in    STD_ULOGIC;
      K                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of JKFF : entity is TRUE;
end JKFF;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library VF1;
architecture VITAL_VF of JKFF is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL J_ipd	 : STD_ULOGIC := 'X';
   SIGNAL K_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL J_CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL K_CLK_dly	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (J_ipd, J, tipd_J);
   VitalWireDelay (K_ipd, K, tipd_K);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   VitalSignalDelay (CLK_dly, CLK_ipd, ticd_CLK);
   VitalSignalDelay (J_CLK_dly, J_ipd, tisd_J_CLK);
   VitalSignalDelay (K_CLK_dly, K_ipd, tisd_K_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (CLK_dly, J_CLK_dly, K_CLK_dly)

   -- timing check results
   VARIABLE Tviol_J_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_J_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_K_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_K_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 4);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_J_CLK_posedge,
          TimingData              => Tmkr_J_CLK_posedge,
          TestSignal              => J_CLK_dly,
          TestSignalName          => "J",
          TestDelay               => tisd_J_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          SetupHigh               => tsetup_J_CLK_noedge_posedge,
          SetupLow                => tsetup_J_CLK_noedge_posedge,
          HoldHigh                => thold_J_CLK_noedge_posedge,
          HoldLow                 => thold_J_CLK_noedge_posedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JKFF",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_K_CLK_posedge,
          TimingData              => Tmkr_K_CLK_posedge,
          TestSignal              => K_CLK_dly,
          TestSignalName          => "K",
          TestDelay               => tisd_K_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          SetupHigh               => tsetup_K_CLK_noedge_posedge,
          SetupLow                => tsetup_K_CLK_noedge_posedge,
          HoldHigh                => thold_K_CLK_noedge_posedge,
          HoldLow                 => thold_K_CLK_noedge_posedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JKFF",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_dly,
          TestSignalName          => "CLK",
          TestDelay               => ticd_CLK,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/JKFF",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_J_CLK_posedge or Tviol_K_CLK_posedge or Pviol_CLK;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => jkfftab,
        DataIn => (
               CLK_dly, J_CLK_dly, K_CLK_dly, '1','1'));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (CLK_dly'last_event, tpd_CLK_Q, TRUE)),
       Mode => VitalInertial,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;

configuration CFG_JKFF_VITAL of JKFF is 
        for VITAL_VF
        end for; 
end CFG_JKFF_VITAL;
----- VITAL model for cell JKFFR -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;

LIBRARY VF1 ;
use VF1.VLOGTOVITAL_TABLES.all;



-- entity declaration --
entity JKFFR is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_R_Q                        :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tsetup_J_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      thold_J_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      tsetup_K_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      thold_K_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      trecovery_R_CLK_posedge_posedge :	VitalDelayType := 2.200 ns;
      thold_R_CLK_posedge_posedge    :	VitalDelayType := 2.200 ns;
      tpw_CLK_posedge         :	VitalDelayType := 4.400 ns;
      tperiod_CLK_posedge             :	VitalDelayType := 8.800 ns;
      ticd_CLK                       :	VitalDelayType := 0.000 ns;
      tisd_J_CLK                     :	VitalDelayType := 0.000 ns;
      tisd_K_CLK                     :	VitalDelayType := 0.000 ns;
      tisd_R_CLK                     :	VitalDelayType := 0.000 ns;
      tipd_J                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_K                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_R                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      J                              :	in    STD_ULOGIC;
      K                              :	in    STD_ULOGIC;
      R                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of JKFFR : entity is TRUE;
end JKFFR;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library VF1;
architecture VITAL_VF of JKFFR is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL J_ipd	 : STD_ULOGIC := 'X';
   SIGNAL K_ipd	 : STD_ULOGIC := 'X';
   SIGNAL R_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL J_CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL K_CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL R_CLK_dly	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (J_ipd, J, tipd_J);
   VitalWireDelay (K_ipd, K, tipd_K);
   VitalWireDelay (R_ipd, R, tipd_R);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   VitalSignalDelay (CLK_dly, CLK_ipd, ticd_CLK);
   VitalSignalDelay (J_CLK_dly, J_ipd, tisd_J_CLK);
   VitalSignalDelay (K_CLK_dly, K_ipd, tisd_K_CLK);
   VitalSignalDelay (R_CLK_dly, R_ipd, tisd_R_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (CLK_dly, J_CLK_dly, K_CLK_dly, R_CLK_dly)

   -- timing check results
   VARIABLE Tviol_J_CLK_R_EQ_1_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_J_CLK_R_EQ_1_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_K_CLK_R_EQ_1_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_K_CLK_R_EQ_1_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_R_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_R_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK_R_EQ_1	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK_R_EQ_1	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 4);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_J_CLK_R_EQ_1_posedge,
          TimingData              => Tmkr_J_CLK_R_EQ_1_posedge,
          TestSignal              => J_CLK_dly,
          TestSignalName          => "J",
          TestDelay               => tisd_J_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          SetupHigh               => tsetup_J_CLK_noedge_posedge,
          SetupLow                => tsetup_J_CLK_noedge_posedge,
          HoldHigh                => thold_J_CLK_noedge_posedge,
          HoldLow                 => thold_J_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(R_CLK_dly) = '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JKFFR",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_K_CLK_R_EQ_1_posedge,
          TimingData              => Tmkr_K_CLK_R_EQ_1_posedge,
          TestSignal              => K_CLK_dly,
          TestSignalName          => "K",
          TestDelay               => tisd_K_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          SetupHigh               => tsetup_K_CLK_noedge_posedge,
          SetupLow                => tsetup_K_CLK_noedge_posedge,
          HoldHigh                => thold_K_CLK_noedge_posedge,
          HoldLow                 => thold_K_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(R_CLK_dly) = '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JKFFR",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_R_CLK_posedge,
          TimingData              => Tmkr_R_CLK_posedge,
          TestSignal              => R_CLK_dly,
          TestSignalName          => "R",
          TestDelay               => tisd_R_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          Recovery                => trecovery_R_CLK_posedge_posedge,
          Removal                 => thold_R_CLK_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JKFFR",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK_R_EQ_1,
          PeriodData              => PInfo_CLK_R_EQ_1,
          TestSignal              => CLK_dly,
          TestSignalName          => "CLK",
          TestDelay               => ticd_CLK,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TO_X01((R_CLK_dly) ) = '1',
          HeaderMsg               => InstancePath & "/JKFFR",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_J_CLK_R_EQ_1_posedge or Tviol_K_CLK_R_EQ_1_posedge or Pviol_CLK_R_EQ_1 or Tviol_R_CLK_posedge;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => jkfftab,
        DataIn => (
               CLK_dly, J_CLK_dly, K_CLK_dly, '1', R_CLK_dly));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (R_CLK_dly'last_event, tpd_R_Q, TRUE),
                 1 => (CLK_dly'last_event, tpd_CLK_Q, TRUE)),
       Mode => VitalInertial,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;

configuration CFG_JKFFR_VITAL of JKFFR is 
        for VITAL_VF
        end for; 
end CFG_JKFFR_VITAL;
----- VITAL model for cell JKFFRH -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;

LIBRARY VF1 ;
use VF1.VLOGTOVITAL_TABLES.all;



-- entity declaration --
entity JKFFRH is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_R_Q                        :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tsetup_J_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      thold_J_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      tsetup_K_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      thold_K_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      trecovery_R_CLK_negedge_posedge :	VitalDelayType := 2.200 ns;
      thold_R_CLK_negedge_posedge    :	VitalDelayType := 2.200 ns;
      tpw_CLK_posedge         :	VitalDelayType := 4.400 ns;
      tpw_R_posedge         :	VitalDelayType := 4.400 ns;
      tperiod_CLK_posedge             :	VitalDelayType := 8.800 ns;
      ticd_CLK                       :	VitalDelayType := 0.000 ns;
      tisd_J_CLK                     :	VitalDelayType := 0.000 ns;
      tisd_K_CLK                     :	VitalDelayType := 0.000 ns;
      tisd_R_CLK                     :	VitalDelayType := 0.000 ns;
      tipd_J                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_K                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_R                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      J                              :	in    STD_ULOGIC;
      K                              :	in    STD_ULOGIC;
      R                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of JKFFRH : entity is TRUE;
end JKFFRH;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library VF1;
architecture VITAL_VF of JKFFRH is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL J_ipd	 : STD_ULOGIC := 'X';
   SIGNAL K_ipd	 : STD_ULOGIC := 'X';
   SIGNAL R_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL J_CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL K_CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL R_CLK_dly	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (J_ipd, J, tipd_J);
   VitalWireDelay (K_ipd, K, tipd_K);
   VitalWireDelay (R_ipd, R, tipd_R);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   VitalSignalDelay (CLK_dly, CLK_ipd, ticd_CLK);
   VitalSignalDelay (J_CLK_dly, J_ipd, tisd_J_CLK);
   VitalSignalDelay (K_CLK_dly, K_ipd, tisd_K_CLK);
   VitalSignalDelay (R_CLK_dly, R_ipd, tisd_R_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (CLK_dly, J_CLK_dly, K_CLK_dly, R_CLK_dly)

   -- timing check results
   VARIABLE Tviol_J_CLK_R_EQ_0_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_J_CLK_R_EQ_0_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_K_CLK_R_EQ_0_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_K_CLK_R_EQ_0_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_R_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_R_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK_R_EQ_0	: STD_ULOGIC := '0';
   VARIABLE Pviol_R	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK_R_EQ_0	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE PInfo_R	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 4);
   VARIABLE R_inverted : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_J_CLK_R_EQ_0_posedge,
          TimingData              => Tmkr_J_CLK_R_EQ_0_posedge,
          TestSignal              => J_CLK_dly,
          TestSignalName          => "J",
          TestDelay               => tisd_J_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          SetupHigh               => tsetup_J_CLK_noedge_posedge,
          SetupLow                => tsetup_J_CLK_noedge_posedge,
          HoldHigh                => thold_J_CLK_noedge_posedge,
          HoldLow                 => thold_J_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(R_CLK_dly) = '0',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JKFFRH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_K_CLK_R_EQ_0_posedge,
          TimingData              => Tmkr_K_CLK_R_EQ_0_posedge,
          TestSignal              => K_CLK_dly,
          TestSignalName          => "K",
          TestDelay               => tisd_K_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          SetupHigh               => tsetup_K_CLK_noedge_posedge,
          SetupLow                => tsetup_K_CLK_noedge_posedge,
          HoldHigh                => thold_K_CLK_noedge_posedge,
          HoldLow                 => thold_K_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(R_CLK_dly) = '0',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JKFFRH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_R_CLK_posedge,
          TimingData              => Tmkr_R_CLK_posedge,
          TestSignal              => R_CLK_dly,
          TestSignalName          => "R",
          TestDelay               => tisd_R_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          Recovery                => trecovery_R_CLK_negedge_posedge,
          Removal                 => thold_R_CLK_negedge_posedge,
          ActiveLow               => FALSE,
          CheckEnabled            => TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JKFFRH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_R,
          PeriodData              => PInfo_R,
          TestSignal              => R_CLK_dly,
          TestSignalName          => "R",
          TestDelay               => tisd_R_CLK,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_R_posedge,
          CheckEnabled            => TRUE, 
          HeaderMsg               => InstancePath & "/JKFFRH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK_R_EQ_0,
          PeriodData              => PInfo_CLK_R_EQ_0,
          TestSignal              => CLK_dly,
          TestSignalName          => "CLK",
          TestDelay               => ticd_CLK,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TO_X01(R_CLK_dly ) = '0',
          HeaderMsg               => InstancePath & "/JKFFRH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_J_CLK_R_EQ_0_posedge or Tviol_R_CLK_posedge or Pviol_CLK_R_EQ_0 or Tviol_K_CLK_R_EQ_0_posedge or Pviol_R;
      R_inverted := (NOT R_CLK_dly);
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => jkfftab,
        DataIn => (
               CLK_dly, J_CLK_dly, K_CLK_dly, '1', R_inverted));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (R_CLK_dly'last_event, tpd_R_Q, TRUE),
                 1 => (CLK_dly'last_event, tpd_CLK_Q, TRUE)),
       Mode => VitalInertial,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;

configuration CFG_JKFFRH_VITAL of JKFFRH is 
        for VITAL_VF
        end for; 
end CFG_JKFFRH_VITAL;
----- VITAL model for cell JKFFRS -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;
LIBRARY VF1 ;
use VF1.VLOGTOVITAL_TABLES.all;


-- entity declaration --
entity JKFFRS is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_R_Q                        :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tpd_S_Q                        :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tsetup_J_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      thold_J_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      tsetup_K_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      thold_K_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      trecovery_R_CLK_posedge_posedge :	VitalDelayType := 2.200 ns;
      thold_R_CLK_posedge_posedge :	VitalDelayType := 2.200 ns;
      trecovery_S_CLK_posedge_posedge :	VitalDelayType := 2.200 ns;
      thold_S_CLK_posedge_posedge :	VitalDelayType := 2.200 ns;
      tpw_CLK_posedge :	VitalDelayType := 4.400 ns;
      tpw_R_negedge :	VitalDelayType := 4.400 ns;
      tpw_S_negedge :	VitalDelayType := 4.400 ns;
      tperiod_CLK_posedge   :	VitalDelayType := 8.800 ns;
      ticd_CLK                       :	VitalDelayType := 0.000 ns;
      tisd_J_CLK                     :	VitalDelayType := 0.000 ns;
      tisd_K_CLK                     :	VitalDelayType := 0.000 ns;
      tisd_R_CLK                     :	VitalDelayType := 0.000 ns;
      tisd_S_CLK                     :	VitalDelayType := 0.000 ns;
      tipd_J                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_K                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_R                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      J                              :	in    STD_ULOGIC;
      K                              :	in    STD_ULOGIC;
      R                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of JKFFRS : entity is TRUE;
end JKFFRS;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library VF1;
use VF1.VLOGTOVITAL_TABLES.all;
architecture VITAL_VF of JKFFRS is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL J_ipd	 : STD_ULOGIC := 'X';
   SIGNAL K_ipd	 : STD_ULOGIC := 'X';
   SIGNAL R_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL J_CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL K_CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL R_CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL S_CLK_dly	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (J_ipd, J, tipd_J);
   VitalWireDelay (K_ipd, K, tipd_K);
   VitalWireDelay (R_ipd, R, tipd_R);
   VitalWireDelay (S_ipd, S, tipd_S);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   VitalSignalDelay (CLK_dly, CLK_ipd, ticd_CLK);
   VitalSignalDelay (J_CLK_dly, J_ipd, tisd_J_CLK);
   VitalSignalDelay (K_CLK_dly, K_ipd, tisd_K_CLK);
   VitalSignalDelay (R_CLK_dly, R_ipd, tisd_R_CLK);
   VitalSignalDelay (S_CLK_dly, S_ipd, tisd_S_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (CLK_dly, J_CLK_dly, K_CLK_dly, R_CLK_dly, S_CLK_dly)

   -- timing check results
   VARIABLE Tviol_J_CLK_R_EQ_1_AN_S_EQ_1_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_J_CLK_R_EQ_1_AN_S_EQ_1_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_K_CLK_R_EQ_1_AN_S_EQ_1_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_K_CLK_R_EQ_1_AN_S_EQ_1_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_R_CLK_S_EQ_1_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_R_CLK_S_EQ_1_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S_CLK_R_EQ_1_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S_CLK_R_EQ_1_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK_R_EQ_1_AN_S_EQ_1	: STD_ULOGIC := '0';
   VARIABLE Pviol_R	: STD_ULOGIC := '0';
   VARIABLE Pviol_S	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK_R_EQ_1_AN_S_EQ_1	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE PInfo_R	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE PInfo_S	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(1 to 5);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_J_CLK_R_EQ_1_AN_S_EQ_1_posedge,
          TimingData              => Tmkr_J_CLK_R_EQ_1_AN_S_EQ_1_posedge,
          TestSignal              => J_CLK_dly,
          TestSignalName          => "J",
          TestDelay               => tisd_J_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          SetupHigh               => tsetup_J_CLK_noedge_posedge,
          SetupLow                => tsetup_J_CLK_noedge_posedge,
          HoldHigh                => thold_J_CLK_noedge_posedge,
          HoldLow                 => thold_J_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((S_CLK_dly) AND (R_CLK_dly)) /= '0',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JKFFRS",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_K_CLK_R_EQ_1_AN_S_EQ_1_posedge,
          TimingData              => Tmkr_K_CLK_R_EQ_1_AN_S_EQ_1_posedge,
          TestSignal              => K_CLK_dly,
          TestSignalName          => "K",
          TestDelay               => tisd_K_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          SetupHigh               => tsetup_K_CLK_noedge_posedge,
          SetupLow                => tsetup_K_CLK_noedge_posedge,
          HoldHigh                => thold_K_CLK_noedge_posedge,
          HoldLow                 => thold_K_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((S_CLK_dly) AND (R_CLK_dly)) /= '0',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JKFFRS",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_R_CLK_S_EQ_1_posedge,
          TimingData              => Tmkr_R_CLK_S_EQ_1_posedge,
          TestSignal              => R_CLK_dly,
          TestSignalName          => "R",
          TestDelay               => tisd_R_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          Recovery                => trecovery_R_CLK_posedge_posedge,
          Removal                 => thold_R_CLK_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TO_X01(S_CLK_dly) /= '0',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JKFFRS",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_S_CLK_R_EQ_1_posedge,
          TimingData              => Tmkr_S_CLK_R_EQ_1_posedge,
          TestSignal              => S_CLK_dly,
          TestSignalName          => "S",
          TestDelay               => tisd_S_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          Recovery                => trecovery_S_CLK_posedge_posedge,
          Removal                 => thold_S_CLK_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TO_X01(R_CLK_dly) /= '0',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JKFFRS",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_S,
          PeriodData              => PInfo_S,
          TestSignal              => S_CLK_dly,
          TestSignalName          => "S",
          TestDelay               => tisd_S_CLK,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_S_negedge,
          CheckEnabled            => TRUE, 
          HeaderMsg               => InstancePath & "/JKFRS",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_R,
          PeriodData              => PInfo_R,
          TestSignal              => R_CLK_dly,
          TestSignalName          => "R",
          TestDelay               => tisd_R_CLK,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_R_negedge,
          CheckEnabled            => TRUE, 
          HeaderMsg               => InstancePath & "/JKRS",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK_R_EQ_1_AN_S_EQ_1,
          PeriodData              => PInfo_CLK_R_EQ_1_AN_S_EQ_1,
          TestSignal              => CLK_dly,
          TestSignalName          => "CLK",
          TestDelay               => ticd_CLK,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TO_X01(( (NOT S_CLK_dly) ) OR ( (NOT R_CLK_dly) )
                            ) /= '1',
          HeaderMsg               => InstancePath & "/JKFFRS",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_J_CLK_R_EQ_1_AN_S_EQ_1_posedge or Tviol_K_CLK_R_EQ_1_AN_S_EQ_1_posedge or Tviol_R_CLK_S_EQ_1_posedge or Pviol_CLK_R_EQ_1_AN_S_EQ_1 or Tviol_S_CLK_R_EQ_1_posedge or Pviol_R or Pviol_S;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => jkfftab,
        DataIn => (
                CLK_dly,J_CLK_dly,K_CLK_dly,S_CLK_dly,R_CLK_dly));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (R_CLK_dly'last_event, tpd_R_Q, TRUE),
                 1 => (S_CLK_dly'last_event, tpd_S_Q, TRUE),
                 2 => (CLK_dly'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;

configuration CFG_JKFFRS_VITAL of JKFFRS is 
        for VITAL_VF
        end for; 
end CFG_JKFFRS_VITAL;
----- VITAL model for cell JKFFRSH -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;
LIBRARY VF1 ;
use VF1.VLOGTOVITAL_TABLES.all;

-- entity declaration --
entity JKFFRSH is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_R_Q                        :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tpd_S_Q                        :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tsetup_J_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      thold_J_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      tsetup_K_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      thold_K_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      trecovery_R_CLK_negedge_posedge :	VitalDelayType := 2.200 ns;
      thold_R_CLK_negedge_posedge :	VitalDelayType := 2.200 ns;
      trecovery_S_CLK_negedge_posedge :	VitalDelayType := 2.200 ns;
      thold_S_CLK_negedge_posedge :	VitalDelayType := 2.200 ns;
      tpw_CLK_posedge :	VitalDelayType := 4.400 ns;
      tpw_R_posedge :	VitalDelayType := 4.400 ns;
      tpw_S_posedge :	VitalDelayType := 4.400 ns;
      tperiod_CLK_posedge   :	VitalDelayType := 8.800 ns;
      ticd_CLK                       :	VitalDelayType := 0.000 ns;
      tisd_J_CLK                     :	VitalDelayType := 0.000 ns;
      tisd_K_CLK                     :	VitalDelayType := 0.000 ns;
      tisd_R_CLK                     :	VitalDelayType := 0.000 ns;
      tisd_S_CLK                     :	VitalDelayType := 0.000 ns;
      tipd_J                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_K                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_R                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      J                              :	in    STD_ULOGIC;
      K                              :	in    STD_ULOGIC;
      R                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of JKFFRSH : entity is TRUE;
end JKFFRSH;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library VF1;
architecture VITAL_VF of JKFFRSH is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL J_ipd	 : STD_ULOGIC := 'X';
   SIGNAL K_ipd	 : STD_ULOGIC := 'X';
   SIGNAL R_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL J_CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL K_CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL R_CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL S_CLK_dly	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (J_ipd, J, tipd_J);
   VitalWireDelay (K_ipd, K, tipd_K);
   VitalWireDelay (R_ipd, R, tipd_R);
   VitalWireDelay (S_ipd, S, tipd_S);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   VitalSignalDelay (CLK_dly, CLK_ipd, ticd_CLK);
   VitalSignalDelay (J_CLK_dly, J_ipd, tisd_J_CLK);
   VitalSignalDelay (K_CLK_dly, K_ipd, tisd_K_CLK);
   VitalSignalDelay (R_CLK_dly, R_ipd, tisd_R_CLK);
   VitalSignalDelay (S_CLK_dly, S_ipd, tisd_S_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (CLK_dly, J_CLK_dly, K_CLK_dly, R_CLK_dly, S_CLK_dly)

   -- timing check results
   VARIABLE Tviol_J_CLK_R_EQ_0_AN_S_EQ_0_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_J_CLK_R_EQ_0_AN_S_EQ_0_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_K_CLK_R_EQ_0_AN_S_EQ_0_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_K_CLK_R_EQ_0_AN_S_EQ_0_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_R_CLK_S_EQ_0_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_R_CLK_S_EQ_0_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S_CLK_R_EQ_0_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S_CLK_R_EQ_0_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK_R_EQ_0_AN_S_EQ_0	: STD_ULOGIC := '0';
   VARIABLE Pviol_R	: STD_ULOGIC := '0';
   VARIABLE Pviol_S	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK_R_EQ_0_AN_S_EQ_0	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE PInfo_R	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE PInfo_S	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(1 to 5);
   VARIABLE J_delayed : STD_ULOGIC := 'X';
   VARIABLE K_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE R_inverted : STD_ULOGIC := 'X';
   VARIABLE S_inverted  : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_J_CLK_R_EQ_0_AN_S_EQ_0_posedge,
          TimingData              => Tmkr_J_CLK_R_EQ_0_AN_S_EQ_0_posedge,
          TestSignal              => J_CLK_dly,
          TestSignalName          => "J",
          TestDelay               => tisd_J_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          SetupHigh               => tsetup_J_CLK_noedge_posedge,
          SetupLow                => tsetup_J_CLK_noedge_posedge,
          HoldHigh                => thold_J_CLK_noedge_posedge,
          HoldLow                 => thold_J_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(((NOT S_CLK_dly)) AND ((NOT R_CLK_dly))) /=
                            '0',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JKFFRSH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_K_CLK_R_EQ_0_AN_S_EQ_0_posedge,
          TimingData              => Tmkr_K_CLK_R_EQ_0_AN_S_EQ_0_posedge,
          TestSignal              => K_CLK_dly,
          TestSignalName          => "K",
          TestDelay               => tisd_K_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          SetupHigh               => tsetup_K_CLK_noedge_posedge,
          SetupLow                => tsetup_K_CLK_noedge_posedge,
          HoldHigh                => thold_K_CLK_noedge_posedge,
          HoldLow                 => thold_K_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(((NOT S_CLK_dly)) AND ((NOT R_CLK_dly))) /=
                            '0',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JKFFRSH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_R_CLK_S_EQ_0_posedge,
          TimingData              => Tmkr_R_CLK_S_EQ_0_posedge,
          TestSignal              => R_CLK_dly,
          TestSignalName          => "R",
          TestDelay               => tisd_R_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          Recovery                => trecovery_R_CLK_negedge_posedge,
          Removal                 => thold_R_CLK_negedge_posedge,
          ActiveLow               => FALSE,
          CheckEnabled            => 
                           TO_X01((NOT S_CLK_dly)) /= '0',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JKFFRSH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_S_CLK_R_EQ_0_posedge,
          TimingData              => Tmkr_S_CLK_R_EQ_0_posedge,
          TestSignal              => S_CLK_dly,
          TestSignalName          => "S",
          TestDelay               => tisd_S_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          Recovery                => trecovery_S_CLK_negedge_posedge,
          Removal                 => thold_S_CLK_negedge_posedge,
          ActiveLow               => FALSE,
          CheckEnabled            => 
                           TO_X01((NOT R_CLK_dly)) /= '0',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JKFFRSH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_S,
          PeriodData              => PInfo_S,
          TestSignal              => S_CLK_dly,
          TestSignalName          => "S",
          TestDelay               => tisd_S_CLK,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_S_posedge,
          CheckEnabled            => TRUE, 
          HeaderMsg               => InstancePath & "/JKFFRSH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_R,
          PeriodData              => PInfo_R,
          TestSignal              => R_CLK_dly,
          TestSignalName          => "R",
          TestDelay               => tisd_R_CLK,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_R_posedge,
          CheckEnabled            => TRUE, 
          HeaderMsg               => InstancePath & "/JKFFRSH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK_R_EQ_0_AN_S_EQ_0,
          PeriodData              => PInfo_CLK_R_EQ_0_AN_S_EQ_0,
          TestSignal              => CLK_dly,
          TestSignalName          => "CLK",
          TestDelay               => ticd_CLK,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TO_X01(( S_CLK_dly ) OR ( R_CLK_dly ) ) /= '1',
          HeaderMsg               => InstancePath & "/JKFFRSH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_J_CLK_R_EQ_0_AN_S_EQ_0_posedge or Tviol_K_CLK_R_EQ_0_AN_S_EQ_0_posedge or Tviol_S_CLK_R_EQ_0_posedge or Pviol_CLK_R_EQ_0_AN_S_EQ_0 or Tviol_R_CLK_S_EQ_0_posedge or Pviol_R or Pviol_S;
      J_delayed := J_CLK_dly;
      K_delayed := K_CLK_dly;
      CLK_delayed := CLK_dly;
      R_inverted :=NOT R_CLK_dly;
      S_inverted :=NOT S_CLK_dly;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => jkfftab,
        DataIn => (
               CLK_dly,J_CLK_dly,K_CLK_dly,S_inverted,R_inverted));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (R_CLK_dly'last_event, tpd_R_Q, TRUE),
                 1 => (S_CLK_dly'last_event, tpd_S_Q, TRUE),
                 2 => (CLK_dly'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;

configuration CFG_JKFFRSH_VITAL of JKFFRSH is 
        for VITAL_VF
        end for; 
end CFG_JKFFRSH_VITAL;
----- VITAL model for cell JKFFRSS -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;

LIBRARY VF1 ;
use VF1.VLOGTOVITAL_TABLES.all;



-- entity declaration --
entity JKFFRSS is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_R_Q                        :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tpd_S_Q                        :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tsetup_J_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      thold_J_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      tsetup_K_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      thold_K_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      trecovery_R_CLK_posedge_posedge :	VitalDelayType := 2.200 ns;
      thold_R_CLK_posedge_posedge :	VitalDelayType := 2.200 ns;
      trecovery_S_CLK_posedge_posedge :	VitalDelayType := 2.200 ns;
      thold_S_CLK_posedge_posedge :	VitalDelayType := 2.200 ns;
      tpw_CLK_posedge :	VitalDelayType := 4.400 ns;
      tperiod_CLK_posedge  :	VitalDelayType := 8.800 ns;
      ticd_CLK                       :	VitalDelayType := 0.000 ns;
      tisd_J_CLK                     :	VitalDelayType := 0.000 ns;
      tisd_K_CLK                     :	VitalDelayType := 0.000 ns;
      tisd_R_CLK                     :	VitalDelayType := 0.000 ns;
      tisd_S_CLK                     :	VitalDelayType := 0.000 ns;
      tipd_J                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_K                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_R                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      J                              :	in    STD_ULOGIC;
      K                              :	in    STD_ULOGIC;
      R                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of JKFFRSS : entity is TRUE;
end JKFFRSS;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library VF1;
architecture VITAL_VF of JKFFRSS is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL J_ipd	 : STD_ULOGIC := 'X';
   SIGNAL K_ipd	 : STD_ULOGIC := 'X';
   SIGNAL R_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL J_CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL K_CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL R_CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL S_CLK_dly	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (J_ipd, J, tipd_J);
   VitalWireDelay (K_ipd, K, tipd_K);
   VitalWireDelay (R_ipd, R, tipd_R);
   VitalWireDelay (S_ipd, S, tipd_S);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   VitalSignalDelay (CLK_dly, CLK_ipd, ticd_CLK);
   VitalSignalDelay (J_CLK_dly, J_ipd, tisd_J_CLK);
   VitalSignalDelay (K_CLK_dly, K_ipd, tisd_K_CLK);
   VitalSignalDelay (R_CLK_dly, R_ipd, tisd_R_CLK);
   VitalSignalDelay (S_CLK_dly, S_ipd, tisd_S_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (CLK_dly, J_CLK_dly, K_CLK_dly, R_CLK_dly, S_CLK_dly)

   -- timing check results
   VARIABLE Tviol_J_CLK_R_EQ_1_ANB_S_EQ_1_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_J_CLK_R_EQ_1_ANB_S_EQ_1_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_K_CLK_R_EQ_1_ANB_S_EQ_1_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_K_CLK_R_EQ_1_ANB_S_EQ_1_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_R_CLK_S_EQ_1_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_R_CLK_S_EQ_1_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S_CLK_R_EQ_1_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S_CLK_R_EQ_1_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK_R_EQ_1_ANB_S_EQ_1	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK_R_EQ_1_ANB_S_EQ_1	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 4);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);
   VARIABLE NOT_S_zd : STD_ULOGIC := '0';
   VARIABLE J_in_zd : STD_ULOGIC := '0';
   VARIABLE K_in_zd : STD_ULOGIC := '0';

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_J_CLK_R_EQ_1_ANB_S_EQ_1_posedge,
          TimingData              => Tmkr_J_CLK_R_EQ_1_ANB_S_EQ_1_posedge,
          TestSignal              => J_CLK_dly,
          TestSignalName          => "J",
          TestDelay               => tisd_J_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          SetupHigh               => tsetup_J_CLK_noedge_posedge,
          SetupLow                => tsetup_J_CLK_noedge_posedge,
          HoldHigh                => thold_J_CLK_noedge_posedge,
          HoldLow                 => thold_J_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((S_CLK_dly) AND (R_CLK_dly)) = '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JKFFRSS",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_K_CLK_R_EQ_1_ANB_S_EQ_1_posedge,
          TimingData              => Tmkr_K_CLK_R_EQ_1_ANB_S_EQ_1_posedge,
          TestSignal              => K_CLK_dly,
          TestSignalName          => "K",
          TestDelay               => tisd_K_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          SetupHigh               => tsetup_K_CLK_noedge_posedge,
          SetupLow                => tsetup_K_CLK_noedge_posedge,
          HoldHigh                => thold_K_CLK_noedge_posedge,
          HoldLow                 => thold_K_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((S_CLK_dly) AND (R_CLK_dly)) = '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JKFFRSS",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_R_CLK_S_EQ_1_posedge,
          TimingData              => Tmkr_R_CLK_S_EQ_1_posedge,
          TestSignal              => R_CLK_dly,
          TestSignalName          => "R",
          TestDelay               => tisd_R_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          Recovery                => trecovery_R_CLK_posedge_posedge,
          Removal                 => thold_R_CLK_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TO_X01(S_CLK_dly) = '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JKFFRSS",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_S_CLK_R_EQ_1_posedge,
          TimingData              => Tmkr_S_CLK_R_EQ_1_posedge,
          TestSignal              => S_CLK_dly,
          TestSignalName          => "S",
          TestDelay               => tisd_S_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          Recovery                => trecovery_S_CLK_posedge_posedge,
          Removal                 => thold_S_CLK_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TO_X01(R_CLK_dly) = '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JKFFRSS",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK_R_EQ_1_ANB_S_EQ_1,
          PeriodData              => PInfo_CLK_R_EQ_1_ANB_S_EQ_1,
          TestSignal              => CLK_dly,
          TestSignalName          => "CLK",
          TestDelay               => ticd_CLK,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TO_X01(( (S_CLK_dly) ) AND ( (R_CLK_dly) )) = '1',
          HeaderMsg               => InstancePath & "/JKFFRSS",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------

        NOT_S_zd := VitalINV (S_CLK_dly);
        J_in_zd := VitalOR2 (NOT_S_zd , J_CLK_dly);
	K_in_zd := VitalAND2 (S_CLK_dly , K_CLK_dly);

      Violation := Tviol_J_CLK_R_EQ_1_ANB_S_EQ_1_posedge or Tviol_K_CLK_R_EQ_1_ANB_S_EQ_1_posedge or Tviol_R_CLK_S_EQ_1_posedge or Tviol_S_CLK_R_EQ_1_posedge or Pviol_CLK_R_EQ_1_ANB_S_EQ_1;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => jkfftab,
        DataIn => (
               CLK_dly, J_in_zd, K_in_zd, '1', R_CLK_dly));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (R_CLK_dly'last_event, tpd_R_Q, TRUE),
                 1 => (S_CLK_dly'last_event, tpd_S_Q, TRUE),
                 2 => (CLK_dly'last_event, tpd_CLK_Q, TRUE)),
       Mode => VitalInertial,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;

configuration CFG_JKFFRSS_VITAL of JKFFRSS is 
        for VITAL_VF
        end for; 
end CFG_JKFFRSS_VITAL;
----- VITAL model for cell JKFFRSSH -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;
LIBRARY VF1 ;
use VF1.VLOGTOVITAL_TABLES.all;



-- entity declaration --
entity JKFFRSSH is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_R_Q                        :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tpd_S_Q                        :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tsetup_J_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      thold_J_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      tsetup_K_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      thold_K_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      trecovery_R_CLK_negedge_posedge :	VitalDelayType := 2.200 ns;
      thold_R_CLK_negedge_posedge :	VitalDelayType := 2.200 ns;
      tsetup_S_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      thold_S_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      tpw_CLK_posedge :	VitalDelayType := 4.400 ns;
      tpw_R_posedge :	VitalDelayType := 4.400 ns;
      tperiod_CLK_posedge  :	VitalDelayType := 8.800 ns;
      ticd_CLK                       :	VitalDelayType := 0.000 ns;
      tisd_J_CLK                     :	VitalDelayType := 0.000 ns;
      tisd_K_CLK                     :	VitalDelayType := 0.000 ns;
      tisd_R_CLK                     :	VitalDelayType := 0.000 ns;
      tisd_S_CLK                     :	VitalDelayType := 0.000 ns;
      tipd_J                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_K                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_R                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      J                              :	in    STD_ULOGIC;
      K                              :	in    STD_ULOGIC;
      R                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of JKFFRSSH : entity is TRUE;
end JKFFRSSH;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library VF1;
architecture VITAL_VF of JKFFRSSH is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL J_ipd	 : STD_ULOGIC := 'X';
   SIGNAL K_ipd	 : STD_ULOGIC := 'X';
   SIGNAL R_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL J_CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL K_CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL R_CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL S_CLK_dly	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (J_ipd, J, tipd_J);
   VitalWireDelay (K_ipd, K, tipd_K);
   VitalWireDelay (R_ipd, R, tipd_R);
   VitalWireDelay (S_ipd, S, tipd_S);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   VitalSignalDelay (CLK_dly, CLK_ipd, ticd_CLK);
   VitalSignalDelay (J_CLK_dly, J_ipd, tisd_J_CLK);
   VitalSignalDelay (K_CLK_dly, K_ipd, tisd_K_CLK);
   VitalSignalDelay (R_CLK_dly, R_ipd, tisd_R_CLK);
   VitalSignalDelay (S_CLK_dly, S_ipd, tisd_S_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (CLK_dly, J_CLK_dly, K_CLK_dly, R_CLK_dly, S_CLK_dly)

   -- timing check results
   VARIABLE Tviol_J_CLK_R_EQ_0_ANB_S_EQ_0_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_J_CLK_R_EQ_0_ANB_S_EQ_0_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_K_CLK_R_EQ_0_ANB_S_EQ_0_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_K_CLK_R_EQ_0_ANB_S_EQ_0_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_R_CLK_S_EQ_0_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_R_CLK_S_EQ_0_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S_CLK_R_EQ_0_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S_CLK_R_EQ_0_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK_R_EQ_0_ANB_S_EQ_0	: STD_ULOGIC := '0';
   VARIABLE Pviol_R	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK_R_EQ_0_ANB_S_EQ_0	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE PInfo_R	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 4);
   VARIABLE R_inverted : STD_ULOGIC := 'X';
   VARIABLE S_inverted : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);
   VARIABLE NOT_S_zd : STD_ULOGIC := '0';
   VARIABLE J_in_zd : STD_ULOGIC := '0';
   VARIABLE K_in_zd : STD_ULOGIC := '0';

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_J_CLK_R_EQ_0_ANB_S_EQ_0_posedge,
          TimingData              => Tmkr_J_CLK_R_EQ_0_ANB_S_EQ_0_posedge,
          TestSignal              => J_CLK_dly,
          TestSignalName          => "J",
          TestDelay               => tisd_J_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          SetupHigh               => tsetup_J_CLK_noedge_posedge,
          SetupLow                => tsetup_J_CLK_noedge_posedge,
          HoldHigh                => thold_J_CLK_noedge_posedge,
          HoldLow                 => thold_J_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(((NOT S_CLK_dly)) AND ((NOT R_CLK_dly))) = '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JKFFRSSH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_K_CLK_R_EQ_0_ANB_S_EQ_0_posedge,
          TimingData              => Tmkr_K_CLK_R_EQ_0_ANB_S_EQ_0_posedge,
          TestSignal              => K_CLK_dly,
          TestSignalName          => "K",
          TestDelay               => tisd_K_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          SetupHigh               => tsetup_K_CLK_noedge_posedge,
          SetupLow                => tsetup_K_CLK_noedge_posedge,
          HoldHigh                => thold_K_CLK_noedge_posedge,
          HoldLow                 => thold_K_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(((NOT S_CLK_dly)) AND ((NOT R_CLK_dly))) = '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JKFFRSSH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_R_CLK_S_EQ_0_posedge,
          TimingData              => Tmkr_R_CLK_S_EQ_0_posedge,
          TestSignal              => R_CLK_dly,
          TestSignalName          => "R",
          TestDelay               => tisd_R_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          Recovery                => trecovery_R_CLK_negedge_posedge,
          Removal                 => thold_R_CLK_negedge_posedge,
          ActiveLow               => FALSE,
          CheckEnabled            => 
                           TO_X01((S_CLK_dly)) = '0',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JKFFRSSH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_S_CLK_R_EQ_0_posedge,
          TimingData              => Tmkr_S_CLK_R_EQ_0_posedge,
          TestSignal              => S_CLK_dly,
          TestSignalName          => "S",
          TestDelay               => tisd_S_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          SetupHigh               => tsetup_S_CLK_noedge_posedge,
          SetupLow                => tsetup_S_CLK_noedge_posedge,
          HoldHigh                => thold_S_CLK_noedge_posedge,
          HoldLow                 => thold_S_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((R_CLK_dly)) = '0',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JKFFRSSH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_R,
          PeriodData              => PInfo_R,
          TestSignal              => R_CLK_dly,
          TestSignalName          => "R",
          TestDelay               => tisd_R_CLK,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_R_posedge,
          CheckEnabled            => TRUE, 
          HeaderMsg               => InstancePath & "/JKFFRSH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK_R_EQ_0_ANB_S_EQ_0,
          PeriodData              => PInfo_CLK_R_EQ_0_ANB_S_EQ_0,
          TestSignal              => CLK_dly,
          TestSignalName          => "CLK",
          TestDelay               => ticd_CLK,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TO_X01(( NOT S_CLK_dly ) AND ( NOT R_CLK_dly ) ) = '1',
          HeaderMsg               => InstancePath & "/JKFFRSSH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------

        NOT_S_zd := VitalINV (S_CLK_dly);
        J_in_zd := VitalOR2 (S_CLK_dly , J_CLK_dly);
        K_in_zd := VitalAND2 (NOT_S_zd , K_CLK_dly);

      Violation := Tviol_J_CLK_R_EQ_0_ANB_S_EQ_0_posedge or Tviol_K_CLK_R_EQ_0_ANB_S_EQ_0_posedge or Tviol_S_CLK_R_EQ_0_posedge or Pviol_CLK_R_EQ_0_ANB_S_EQ_0 or Tviol_R_CLK_S_EQ_0_posedge or Pviol_R;
      R_inverted := (NOT R_CLK_dly);
      S_inverted := (NOT S_CLK_dly);
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => jkfftab,
        DataIn => (
               CLK_dly, J_in_zd, K_in_zd, '1', R_inverted));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (R_CLK_dly'last_event, tpd_R_Q, TRUE),
                 1 => (S_CLK_dly'last_event, tpd_S_Q, TRUE),
                 2 => (CLK_dly'last_event, tpd_CLK_Q, TRUE)),
       Mode => VitalInertial,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;

configuration CFG_JKFFRSSH_VITAL of JKFFRSSH is 
        for VITAL_VF
        end for; 
end CFG_JKFFRSSH_VITAL;
----- VITAL model for cell JKFFS -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;

LIBRARY VF1 ;
use VF1.VLOGTOVITAL_TABLES.all;



-- entity declaration --
entity JKFFS is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_S_Q                        :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tsetup_J_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      thold_J_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      tsetup_K_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      thold_K_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      trecovery_S_CLK_posedge_posedge :	VitalDelayType := 2.200 ns;
      thold_S_CLK_posedge_posedge    :	VitalDelayType := 2.200 ns;
      tpw_CLK_posedge         :	VitalDelayType := 4.400 ns;
      tperiod_CLK_posedge             :	VitalDelayType := 8.800 ns;
      ticd_CLK                       :	VitalDelayType := 0.000 ns;
      tisd_J_CLK                     :	VitalDelayType := 0.000 ns;
      tisd_K_CLK                     :	VitalDelayType := 0.000 ns;
      tisd_S_CLK                     :	VitalDelayType := 0.000 ns;
      tipd_J                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_K                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      J                              :	in    STD_ULOGIC;
      K                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of JKFFS : entity is TRUE;
end JKFFS;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library VF1;
architecture VITAL_VF of JKFFS is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL J_ipd	 : STD_ULOGIC := 'X';
   SIGNAL K_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL J_CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL K_CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL S_CLK_dly	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (J_ipd, J, tipd_J);
   VitalWireDelay (K_ipd, K, tipd_K);
   VitalWireDelay (S_ipd, S, tipd_S);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   VitalSignalDelay (CLK_dly, CLK_ipd, ticd_CLK);
   VitalSignalDelay (J_CLK_dly, J_ipd, tisd_J_CLK);
   VitalSignalDelay (K_CLK_dly, K_ipd, tisd_K_CLK);
   VitalSignalDelay (S_CLK_dly, S_ipd, tisd_S_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (CLK_dly, J_CLK_dly, K_CLK_dly, S_CLK_dly)

   -- timing check results
   VARIABLE Tviol_J_CLK_S_EQ_1_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_J_CLK_S_EQ_1_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_K_CLK_S_EQ_1_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_K_CLK_S_EQ_1_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK_S_EQ_1	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK_S_EQ_1	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 4);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_J_CLK_S_EQ_1_posedge,
          TimingData              => Tmkr_J_CLK_S_EQ_1_posedge,
          TestSignal              => J_CLK_dly,
          TestSignalName          => "J",
          TestDelay               => tisd_J_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          SetupHigh               => tsetup_J_CLK_noedge_posedge,
          SetupLow                => tsetup_J_CLK_noedge_posedge,
          HoldHigh                => thold_J_CLK_noedge_posedge,
          HoldLow                 => thold_J_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(S_CLK_dly) = '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JKFFS",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_K_CLK_S_EQ_1_posedge,
          TimingData              => Tmkr_K_CLK_S_EQ_1_posedge,
          TestSignal              => K_CLK_dly,
          TestSignalName          => "K",
          TestDelay               => tisd_K_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          SetupHigh               => tsetup_K_CLK_noedge_posedge,
          SetupLow                => tsetup_K_CLK_noedge_posedge,
          HoldHigh                => thold_K_CLK_noedge_posedge,
          HoldLow                 => thold_K_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(S_CLK_dly) = '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JKFFS",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_S_CLK_posedge,
          TimingData              => Tmkr_S_CLK_posedge,
          TestSignal              => S_CLK_dly,
          TestSignalName          => "S",
          TestDelay               => tisd_S_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          Recovery                => trecovery_S_CLK_posedge_posedge,
          Removal                 => thold_S_CLK_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JKFFS",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK_S_EQ_1,
          PeriodData              => PInfo_CLK_S_EQ_1,
          TestSignal              => CLK_dly,
          TestSignalName          => "CLK",
          TestDelay               => ticd_CLK,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TO_X01((S_CLK_dly) ) = '1',
          HeaderMsg               => InstancePath & "/JKFFS",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_J_CLK_S_EQ_1_posedge or Tviol_K_CLK_S_EQ_1_posedge or Tviol_S_CLK_posedge or Pviol_CLK_S_EQ_1;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => jkfftab,
        DataIn => (
               CLK_dly, J_CLK_dly, K_CLK_dly, S_CLK_dly, '1'));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (S_CLK_dly'last_event, tpd_S_Q, TRUE),
                 1 => (CLK_dly'last_event, tpd_CLK_Q, TRUE)),
       Mode => VitalInertial,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;

configuration CFG_JKFFS_VITAL of JKFFS is 
        for VITAL_VF
        end for; 
end CFG_JKFFS_VITAL;
----- VITAL model for cell JKFFSH -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;

LIBRARY VF1 ;
use VF1.VLOGTOVITAL_TABLES.all;



-- entity declaration --
entity JKFFSH is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_S_Q                        :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tsetup_J_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      thold_J_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      tsetup_K_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      thold_K_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      trecovery_S_CLK_negedge_posedge :	VitalDelayType := 2.200 ns;
      thold_S_CLK_negedge_posedge    :	VitalDelayType := 2.200 ns;
      tpw_CLK_posedge         :	VitalDelayType := 4.400 ns;
      tpw_S_posedge         :	VitalDelayType := 4.400 ns;
      tperiod_CLK_posedge             :	VitalDelayType := 8.800 ns;
      ticd_CLK                       :	VitalDelayType := 0.000 ns;
      tisd_J_CLK                     :	VitalDelayType := 0.000 ns;
      tisd_K_CLK                     :	VitalDelayType := 0.000 ns;
      tisd_S_CLK                     :	VitalDelayType := 0.000 ns;
      tipd_J                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_K                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      J                              :	in    STD_ULOGIC;
      K                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of JKFFSH : entity is TRUE;
end JKFFSH;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library VF1;
architecture VITAL_VF of JKFFSH is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL J_ipd	 : STD_ULOGIC := 'X';
   SIGNAL K_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL J_CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL K_CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL S_CLK_dly	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (J_ipd, J, tipd_J);
   VitalWireDelay (K_ipd, K, tipd_K);
   VitalWireDelay (S_ipd, S, tipd_S);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   VitalSignalDelay (CLK_dly, CLK_ipd, ticd_CLK);
   VitalSignalDelay (J_CLK_dly, J_ipd, tisd_J_CLK);
   VitalSignalDelay (K_CLK_dly, K_ipd, tisd_K_CLK);
   VitalSignalDelay (S_CLK_dly, S_ipd, tisd_S_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (CLK_dly, J_CLK_dly, K_CLK_dly, S_CLK_dly)

   -- timing check results
   VARIABLE Tviol_J_CLK_S_EQ_0_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_J_CLK_S_EQ_0_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_K_CLK_S_EQ_0_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_K_CLK_S_EQ_0_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK_S_EQ_0	: STD_ULOGIC := '0';
   VARIABLE Pviol_S	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK_S_EQ_0	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE PInfo_S	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 4);
   VARIABLE S_inverted : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_J_CLK_S_EQ_0_posedge,
          TimingData              => Tmkr_J_CLK_S_EQ_0_posedge,
          TestSignal              => J_CLK_dly,
          TestSignalName          => "J",
          TestDelay               => tisd_J_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          SetupHigh               => tsetup_J_CLK_noedge_posedge,
          SetupLow                => tsetup_J_CLK_noedge_posedge,
          HoldHigh                => thold_J_CLK_noedge_posedge,
          HoldLow                 => thold_J_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(S_CLK_dly) = '0',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JKFFSH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_K_CLK_S_EQ_0_posedge,
          TimingData              => Tmkr_K_CLK_S_EQ_0_posedge,
          TestSignal              => K_CLK_dly,
          TestSignalName          => "K",
          TestDelay               => tisd_K_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          SetupHigh               => tsetup_K_CLK_noedge_posedge,
          SetupLow                => tsetup_K_CLK_noedge_posedge,
          HoldHigh                => thold_K_CLK_noedge_posedge,
          HoldLow                 => thold_K_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(S_CLK_dly) = '0',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JKFFSH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_S_CLK_posedge,
          TimingData              => Tmkr_S_CLK_posedge,
          TestSignal              => S_CLK_dly,
          TestSignalName          => "S",
          TestDelay               => tisd_S_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          Recovery                => trecovery_S_CLK_negedge_posedge,
          Removal                 => thold_S_CLK_negedge_posedge,
          ActiveLow               => FALSE,
          CheckEnabled            => TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JKFFSH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_S,
          PeriodData              => PInfo_S,
          TestSignal              => S_CLK_dly,
          TestSignalName          => "S",
          TestDelay               => tisd_S_CLK,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_S_posedge,
          CheckEnabled            => TRUE, 
          HeaderMsg               => InstancePath & "/JKFFSH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK_S_EQ_0,
          PeriodData              => PInfo_CLK_S_EQ_0,
          TestSignal              => CLK_dly,
          TestSignalName          => "CLK",
          TestDelay               => ticd_CLK,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TO_X01(S_CLK_dly ) = '0',
          HeaderMsg               => InstancePath & "/JKFFSH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_J_CLK_S_EQ_0_posedge or Tviol_S_CLK_posedge or Pviol_CLK_S_EQ_0 or Tviol_K_CLK_S_EQ_0_posedge or Pviol_S;
      S_inverted := (NOT S_CLK_dly);
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => jkfftab,
        DataIn => (
               CLK_dly, J_CLK_dly, K_CLK_dly, S_inverted, '1'));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (S_CLK_dly'last_event, tpd_S_Q, TRUE),
                 1 => (CLK_dly'last_event, tpd_CLK_Q, TRUE)),
       Mode => VitalInertial,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;

configuration CFG_JKFFSH_VITAL of JKFFSH is 
        for VITAL_VF
        end for; 
end CFG_JKFFSH_VITAL;
----- VITAL model for cell JTAG -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity JTAG is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tipd_TDI                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_TCLK                      :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_TMOD                      :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      TDI                             :	in    STD_ULOGIC;
      TCLK                           :	in    STD_ULOGIC;
      TMOD                           :	in    STD_ULOGIC;
      TDO                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of JTAG : entity is TRUE;
end JTAG;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library VF1;
architecture VITAL_VF of JTAG is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL TDI_ipd	 : STD_ULOGIC := 'X';
   SIGNAL TCLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL TMOD_ipd	 : STD_ULOGIC := 'X';
   SIGNAL TEMP		 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (TDI_ipd, TDI, tipd_TDI);
   VitalWireDelay (TCLK_ipd, TCLK, tipd_TCLK);
   VitalWireDelay (TMOD_ipd, TMOD, tipd_TMOD);
   end block;

Inst1: VitalIDENT (TDO,TEMP);

end VITAL_VF;

configuration CFG_JTAG_VITAL of JTAG is 
        for VITAL_VF
        end for; 
end CFG_JTAG_VITAL;
----- VITAL model for cell LI -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;

LIBRARY VF1 ;
use VF1.VLOGTOVITAL_TABLES.all;


-- entity declaration --
entity LI is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_D_Q                        :	VitalDelayType01 := (1.230 ns, 1.230 ns);
      tpd_LAT_Q                      :	VitalDelayType01 := (1.230 ns, 1.230 ns);
      tsetup_D_LAT_noedge_negedge    :	VitalDelayType := 0.000 ns;
      thold_D_LAT_noedge_negedge     :	VitalDelayType := 0.530 ns;
      tperiod_LAT_posedge            :	VitalDelayType := 1.320 ns;
      tpw_LAT_posedge                :	VitalDelayType := 0.660 ns;
      ticd_LAT                       :	VitalDelayType := 0.000 ns;
      tisd_D_LAT                     :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_LAT                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      LAT                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of LI : entity is TRUE;
end LI;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library VF1;
architecture VITAL_VF of LI is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL LAT_ipd	 : STD_ULOGIC := 'X';
   SIGNAL LAT_dly	 : STD_ULOGIC := 'X';
   SIGNAL D_LAT_dly	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (LAT_ipd, LAT, tipd_LAT);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   VitalSignalDelay (LAT_dly, LAT_ipd, ticd_LAT);
   VitalSignalDelay (D_LAT_dly, D_ipd, tisd_D_LAT);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (LAT_dly, D_LAT_dly)

   -- timing check results
   VARIABLE Tviol_D_LAT_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_LAT_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_LAT	: STD_ULOGIC := '0';
   VARIABLE PInfo_LAT	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 3);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_LAT_negedge,
          TimingData              => Tmkr_D_LAT_negedge,
          TestSignal              => D_LAT_dly,
          TestSignalName          => "D",
          TestDelay               => tisd_D_LAT,
          RefSignal               => LAT_dly,
          RefSignalName          => "LAT",
          RefDelay                => ticd_LAT,
          SetupHigh               => tsetup_D_LAT_noedge_negedge,
          SetupLow                => tsetup_D_LAT_noedge_negedge,
          HoldHigh                => thold_D_LAT_noedge_negedge,
          HoldLow                 => thold_D_LAT_noedge_negedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/LI",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_LAT,
          PeriodData              => PInfo_LAT,
          TestSignal              => LAT_dly,
          TestSignalName          => "LAT",
          TestDelay               => ticd_LAT,
          Period                  => tperiod_LAT_posedge,
          PulseWidthHigh          => tpw_LAT_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/LI",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_LAT_negedge or Pviol_LAT;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => latchtab,
        DataIn => (
               D_LAT_dly, LAT_dly,'1','1'));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (D_LAT_dly'last_event, tpd_D_Q, TRUE),
                 1 => (LAT_dly'last_event, tpd_LAT_Q, TRUE)),
       Mode => VitalInertial,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;

configuration CFG_LI_VITAL of LI is 
        for VITAL_VF
        end for; 
end CFG_LI_VITAL;
----- VITAL model for cell LIR -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;

LIBRARY VF1 ;
use VF1.VLOGTOVITAL_TABLES.all;



-- entity declaration --
entity LIR is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_D_Q                        :	VitalDelayType01 := (1.230 ns, 1.230 ns);
      tpd_LAT_Q                      :	VitalDelayType01 := (1.230 ns, 1.230 ns);
      tpd_R_Q                        :	VitalDelayType01 := (1.230 ns, 1.230 ns);
      tsetup_D_LAT_noedge_negedge :	VitalDelayType := 0.000 ns;---0.330 ns;
      thold_D_LAT_noedge_negedge :	VitalDelayType := 0.530 ns;
      tpw_LAT_posedge         :	VitalDelayType := 0.660 ns;
      tperiod_LAT_posedge             :	VitalDelayType := 1.320 ns;
      trecovery_R_LAT_posedge_negedge :	VitalDelayType := 0.000 ns;---0.330 ns;
      thold_R_LAT_posedge_negedge    :	VitalDelayType := 0.530 ns;
      ticd_LAT                       :	VitalDelayType := 0.000 ns;
      tisd_D_LAT                     :	VitalDelayType := 0.000 ns;
      tisd_R_LAT                     :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_LAT                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_R                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      LAT                            :	in    STD_ULOGIC;
      R                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of LIR : entity is TRUE;
end LIR;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library VF1;
architecture VITAL_VF of LIR is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL LAT_ipd	 : STD_ULOGIC := 'X';
   SIGNAL R_ipd	 : STD_ULOGIC := 'X';
   SIGNAL LAT_dly	 : STD_ULOGIC := 'X';
   SIGNAL D_LAT_dly	 : STD_ULOGIC := 'X';
   SIGNAL R_LAT_dly	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (LAT_ipd, LAT, tipd_LAT);
   VitalWireDelay (R_ipd, R, tipd_R);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   VitalSignalDelay (LAT_dly, LAT_ipd, ticd_LAT);
   VitalSignalDelay (D_LAT_dly, D_ipd, tisd_D_LAT);
   VitalSignalDelay (R_LAT_dly, R_ipd, tisd_R_LAT);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (LAT_dly, D_LAT_dly, R_LAT_dly)

   -- timing check results
   VARIABLE Tviol_D_LAT_R_EQ_1_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_LAT_R_EQ_1_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_R_LAT_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_R_LAT_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_LAT_R_EQ_1	: STD_ULOGIC := '0';
   VARIABLE PInfo_LAT_R_EQ_1	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 3);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_LAT_R_EQ_1_negedge,
          TimingData              => Tmkr_D_LAT_R_EQ_1_negedge,
          TestSignal              => D_LAT_dly,
          TestSignalName          => "D",
          TestDelay               => tisd_D_LAT,
          RefSignal               => LAT_dly,
          RefSignalName          => "LAT",
          RefDelay                => ticd_LAT,
          SetupHigh               => tsetup_D_LAT_noedge_negedge,
          SetupLow                => tsetup_D_LAT_noedge_negedge,
          HoldHigh                => thold_D_LAT_noedge_negedge,
          HoldLow                 => thold_D_LAT_noedge_negedge,
          CheckEnabled            => 
                           TO_X01(R_LAT_dly) = '0',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/LIR",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_R_LAT_negedge,
          TimingData              => Tmkr_R_LAT_negedge,
          TestSignal              => R_LAT_dly,
          TestSignalName          => "R",
          TestDelay               => tisd_R_LAT,
          RefSignal               => LAT_dly,
          RefSignalName          => "LAT",
          RefDelay                => ticd_LAT,
          Recovery                => trecovery_R_LAT_posedge_negedge,
          Removal                 => thold_R_LAT_posedge_negedge,
          ActiveLow               => TRUE,
          CheckEnabled            => TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/LIR",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_LAT_R_EQ_1,
          PeriodData              => PInfo_LAT_R_EQ_1,
          TestSignal              => LAT_dly,
          TestSignalName          => "LAT",
          TestDelay               => ticd_LAT,
          Period                  => tperiod_LAT_posedge,
          PulseWidthHigh          => tpw_LAT_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TO_X01(R_LAT_dly ) = '0',
          HeaderMsg               => InstancePath & "/LIR",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_LAT_R_EQ_1_negedge or Tviol_R_LAT_negedge or Pviol_LAT_R_EQ_1;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => latchtab,
        DataIn => (
               D_LAT_dly, LAT_dly, NOT(R_LAT_dly),'1'));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (D_LAT_dly'last_event, tpd_D_Q, TRUE),
                 1 => (LAT_dly'last_event, tpd_LAT_Q, TRUE),
                 2 => (R_LAT_dly'last_event, tpd_R_Q, TRUE)),
       Mode => VitalInertial,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;

configuration CFG_LIR_VITAL of LIR is 
        for VITAL_VF
        end for; 
end CFG_LIR_VITAL;
----- VITAL model for cell LIS -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;

LIBRARY VF1 ;
use VF1.VLOGTOVITAL_TABLES.all;



-- entity declaration --
entity LIS is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_D_Q                        :	VitalDelayType01 := (1.230 ns, 1.230 ns);
      tpd_LAT_Q                      :	VitalDelayType01 := (1.230 ns, 1.230 ns);
      tpd_S_Q                        :	VitalDelayType01 := (1.230 ns, 1.230 ns);
      tsetup_D_LAT_noedge_negedge :	VitalDelayType := 0.000 ns;---0.330 ns;
      thold_D_LAT_noedge_negedge :	VitalDelayType := 0.530 ns;
      tpw_LAT_posedge         :	VitalDelayType := 0.660 ns;
      tperiod_LAT_posedge             :	VitalDelayType := 1.320 ns;
      trecovery_S_LAT_posedge_negedge :	VitalDelayType := 0.000 ns;---0.330 ns;
      thold_S_LAT_posedge_negedge    :	VitalDelayType := 0.530 ns;
      ticd_LAT                       :	VitalDelayType := 0.000 ns;
      tisd_D_LAT                     :	VitalDelayType := 0.000 ns;
      tisd_S_LAT                     :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_LAT                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      LAT                            :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of LIS : entity is TRUE;
end LIS;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library VF1;
architecture VITAL_VF of LIS is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL LAT_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S_ipd	 : STD_ULOGIC := 'X';
   SIGNAL LAT_dly	 : STD_ULOGIC := 'X';
   SIGNAL D_LAT_dly	 : STD_ULOGIC := 'X';
   SIGNAL S_LAT_dly	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (LAT_ipd, LAT, tipd_LAT);
   VitalWireDelay (S_ipd, S, tipd_S);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   VitalSignalDelay (LAT_dly, LAT_ipd, ticd_LAT);
   VitalSignalDelay (D_LAT_dly, D_ipd, tisd_D_LAT);
   VitalSignalDelay (S_LAT_dly, S_ipd, tisd_S_LAT);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (LAT_dly, D_LAT_dly, S_LAT_dly)

   -- timing check results
   VARIABLE Tviol_D_LAT_S_EQ_1_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_LAT_S_EQ_1_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S_LAT_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S_LAT_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_LAT_S_EQ_1	: STD_ULOGIC := '0';
   VARIABLE PInfo_LAT_S_EQ_1	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 3);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_LAT_S_EQ_1_negedge,
          TimingData              => Tmkr_D_LAT_S_EQ_1_negedge,
          TestSignal              => D_LAT_dly,
          TestSignalName          => "D",
          TestDelay               => tisd_D_LAT,
          RefSignal               => LAT_dly,
          RefSignalName          => "LAT",
          RefDelay                => ticd_LAT,
          SetupHigh               => tsetup_D_LAT_noedge_negedge,
          SetupLow                => tsetup_D_LAT_noedge_negedge,
          HoldHigh                => thold_D_LAT_noedge_negedge,
          HoldLow                 => thold_D_LAT_noedge_negedge,
          CheckEnabled            => 
                           TO_X01(S_LAT_dly) = '0',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/LIS",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_S_LAT_negedge,
          TimingData              => Tmkr_S_LAT_negedge,
          TestSignal              => S_LAT_dly,
          TestSignalName          => "S",
          TestDelay               => tisd_S_LAT,
          RefSignal               => LAT_dly,
          RefSignalName          => "LAT",
          RefDelay                => ticd_LAT,
          Recovery                => trecovery_S_LAT_posedge_negedge,
          Removal                 => thold_S_LAT_posedge_negedge,
          ActiveLow               => TRUE,
          CheckEnabled            => TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/LIS",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_LAT_S_EQ_1,
          PeriodData              => PInfo_LAT_S_EQ_1,
          TestSignal              => LAT_dly,
          TestSignalName          => "LAT",
          TestDelay               => ticd_LAT,
          Period                  => tperiod_LAT_posedge,
          PulseWidthHigh          => tpw_LAT_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TO_X01(S_LAT_dly ) = '0',
          HeaderMsg               => InstancePath & "/LIS",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_LAT_S_EQ_1_negedge or Tviol_S_LAT_negedge or Pviol_LAT_S_EQ_1;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => latchtab,
        DataIn => (
               D_LAT_dly, LAT_dly, '1',NOT(S_LAT_dly)));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (D_LAT_dly'last_event, tpd_D_Q, TRUE),
                 1 => (LAT_dly'last_event, tpd_LAT_Q, TRUE),
                 2 => (S_LAT_dly'last_event, tpd_S_Q, TRUE)),
       Mode => VitalInertial,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;

configuration CFG_LIS_VITAL of LIS is 
        for VITAL_VF
        end for; 
end CFG_LIS_VITAL;
----- VITAL model for cell MAJOR3 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity MAJOR3 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_I0_O                       :	VitalDelayType01 := (1.250 ns, 1.250 ns);
      tpd_I1_O                       :	VitalDelayType01 := (1.250 ns, 1.250 ns);
      tpd_I2_O                       :	VitalDelayType01 := (1.250 ns, 1.250 ns);
      tipd_I0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I2                        :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      I0                             :	in    STD_ULOGIC;
      I1                             :	in    STD_ULOGIC;
      I2                             :	in    STD_ULOGIC;
      O                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of MAJOR3 : entity is TRUE;
end MAJOR3;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_VF of MAJOR3 is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL I0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I1_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I2_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (I0_ipd, I0, tipd_I0);
   VitalWireDelay (I1_ipd, I1, tipd_I1);
   VitalWireDelay (I2_ipd, I2, tipd_I2);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (I0_ipd, I1_ipd, I2_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS O_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE O_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      O_zd :=
       ((I2_ipd) AND (I1_ipd)) OR ((I1_ipd) AND (I0_ipd)) OR ((I0_ipd) AND
         (I2_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => O,
       GlitchData => O_GlitchData,
       OutSignalName => "O",
       OutTemp => O_zd,
       Paths => (0 => (I0_ipd'last_event, tpd_I0_O, TRUE),
                 1 => (I1_ipd'last_event, tpd_I1_O, TRUE),
                 2 => (I2_ipd'last_event, tpd_I2_O, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;

configuration CFG_MAJOR3_VITAL of MAJOR3 is 
        for VITAL_VF
        end for; 
end CFG_MAJOR3_VITAL;
----- VITAL model for cell MUX2 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity MUX2 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_I0_O                       :	VitalDelayType01 := (1.25 ns, 1.25 ns);
      tpd_I1_O                       :	VitalDelayType01 := (1.25 ns, 1.25 ns);
      tpd_S0_O                      :	VitalDelayType01 := (1.25 ns, 1.25 ns);
      tipd_I0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S0                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      I0                             :	in    STD_ULOGIC;
      I1                             :	in    STD_ULOGIC;
      S0                            :	in    STD_ULOGIC;
      O                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of MUX2 : entity is TRUE;
end MUX2;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library VF1;
architecture VITAL_VF of MUX2 is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL I0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I1_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S0_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (I0_ipd, I0, tipd_I0);
   VitalWireDelay (I1_ipd, I1, tipd_I1);
   VitalWireDelay (S0_ipd, S0, tipd_S0);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (I0_ipd, I1_ipd, S0_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS O_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE O_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      O_zd := VitalMUX
                 (data => (I1_ipd, I0_ipd),
                  dselect => (0 => S0_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => O,
       GlitchData => O_GlitchData,
       OutSignalName => "O",
       OutTemp => O_zd,
       Paths => (0 => (I0_ipd'last_event, tpd_I0_O, TRUE),
                 1 => (I1_ipd'last_event, tpd_I1_O, TRUE),
                 2 => (S0_ipd'last_event, tpd_S0_O, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;

configuration CFG_MUX2_VITAL of MUX2 is 
        for VITAL_VF
        end for; 
end CFG_MUX2_VITAL;
----- VITAL model for cell MUX4 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity MUX4 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_I0_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I1_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I2_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I3_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_S0_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_S1_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tipd_I0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I2                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I3                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      I0                             :	in    STD_ULOGIC;
      I1                             :	in    STD_ULOGIC;
      I2                             :	in    STD_ULOGIC;
      I3                             :	in    STD_ULOGIC;
      S0                             :	in    STD_ULOGIC;
      S1                             :	in    STD_ULOGIC;
      O                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of MUX4 : entity is TRUE;
end MUX4;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library VF1;
architecture VITAL_VF of MUX4 is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL I0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I1_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I2_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I3_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S1_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (I0_ipd, I0, tipd_I0);
   VitalWireDelay (I1_ipd, I1, tipd_I1);
   VitalWireDelay (I2_ipd, I2, tipd_I2);
   VitalWireDelay (I3_ipd, I3, tipd_I3);
   VitalWireDelay (S0_ipd, S0, tipd_S0);
   VitalWireDelay (S1_ipd, S1, tipd_S1);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (I0_ipd, I1_ipd, I2_ipd, I3_ipd, S0_ipd, S1_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS O_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE O_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      O_zd := VitalMUX
                 (data => (I3_ipd, I1_ipd, I2_ipd, I0_ipd),
                  dselect => (S0_ipd, S1_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => O,
       GlitchData => O_GlitchData,
       OutSignalName => "O",
       OutTemp => O_zd,
       Paths => (0 => (I0_ipd'last_event, tpd_I0_O, TRUE),
                 1 => (I1_ipd'last_event, tpd_I1_O, TRUE),
                 2 => (I2_ipd'last_event, tpd_I2_O, TRUE),
                 3 => (I3_ipd'last_event, tpd_I3_O, TRUE),
                 4 => (S0_ipd'last_event, tpd_S0_O, TRUE),
                 5 => (S1_ipd'last_event, tpd_S1_O, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;

configuration CFG_MUX4_VITAL of MUX4 is 
        for VITAL_VF
        end for; 
end CFG_MUX4_VITAL;
----- VITAL model for cell NAN2 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity NAN2 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_I0_O                       :	VitalDelayType01 := (1.25 ns, 1.25 ns);
      tpd_I1_O                       :	VitalDelayType01 := (1.25 ns, 1.25 ns);
      tipd_I0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      I0                             :	in    STD_ULOGIC;
      I1                             :	in    STD_ULOGIC;
      O                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of NAN2 : entity is TRUE;
end NAN2;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library VF1;
architecture VITAL_VF of NAN2 is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL I0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I1_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (I0_ipd, I0, tipd_I0);
   VitalWireDelay (I1_ipd, I1, tipd_I1);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (I0_ipd, I1_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS O_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE O_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      O_zd := ((NOT I1_ipd)) OR ((NOT I0_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => O,
       GlitchData => O_GlitchData,
       OutSignalName => "O",
       OutTemp => O_zd,
       Paths => (0 => (I0_ipd'last_event, tpd_I0_O, TRUE),
                 1 => (I1_ipd'last_event, tpd_I1_O, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;

configuration CFG_NAN2_VITAL of NAN2 is 
        for VITAL_VF
        end for; 
end CFG_NAN2_VITAL;
----- VITAL model for cell NAN3 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity NAN3 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_I0_O                       :	VitalDelayType01 := (1.25 ns, 1.25 ns);
      tpd_I1_O                       :	VitalDelayType01 := (1.25 ns, 1.25 ns);
      tpd_I2_O                       :	VitalDelayType01 := (1.25 ns, 1.25 ns);
      tipd_I0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I2                        :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      I0                             :	in    STD_ULOGIC;
      I1                             :	in    STD_ULOGIC;
      I2                             :	in    STD_ULOGIC;
      O                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of NAN3 : entity is TRUE;
end NAN3;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library VF1;
architecture VITAL_VF of NAN3 is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL I0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I1_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I2_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (I0_ipd, I0, tipd_I0);
   VitalWireDelay (I1_ipd, I1, tipd_I1);
   VitalWireDelay (I2_ipd, I2, tipd_I2);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (I0_ipd, I1_ipd, I2_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS O_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE O_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      O_zd := ((NOT I1_ipd)) OR ((NOT I0_ipd)) OR ((NOT I2_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => O,
       GlitchData => O_GlitchData,
       OutSignalName => "O",
       OutTemp => O_zd,
       Paths => (0 => (I0_ipd'last_event, tpd_I0_O, TRUE),
                 1 => (I1_ipd'last_event, tpd_I1_O, TRUE),
                 2 => (I2_ipd'last_event, tpd_I2_O, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;

configuration CFG_NAN3_VITAL of NAN3 is 
        for VITAL_VF
        end for; 
end CFG_NAN3_VITAL;
----- VITAL model for cell NAN4 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity NAN4 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_I0_O                       :	VitalDelayType01 := (1.80 ns, 1.80 ns);
      tpd_I1_O                       :	VitalDelayType01 := (1.80 ns, 1.80 ns);
      tpd_I2_O                       :	VitalDelayType01 := (1.80 ns, 1.80 ns);
      tpd_I3_O                       :	VitalDelayType01 := (1.80 ns, 1.80 ns);
      tipd_I0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I2                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I3                        :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      I0                             :	in    STD_ULOGIC;
      I1                             :	in    STD_ULOGIC;
      I2                             :	in    STD_ULOGIC;
      I3                             :	in    STD_ULOGIC;
      O                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of NAN4 : entity is TRUE;
end NAN4;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library VF1;
architecture VITAL_VF of NAN4 is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL I0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I1_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I2_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I3_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (I0_ipd, I0, tipd_I0);
   VitalWireDelay (I1_ipd, I1, tipd_I1);
   VitalWireDelay (I2_ipd, I2, tipd_I2);
   VitalWireDelay (I3_ipd, I3, tipd_I3);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (I0_ipd, I1_ipd, I2_ipd, I3_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS O_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE O_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      O_zd :=
       ((NOT I1_ipd)) OR ((NOT I0_ipd)) OR ((NOT I2_ipd)) OR ((NOT I3_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => O,
       GlitchData => O_GlitchData,
       OutSignalName => "O",
       OutTemp => O_zd,
       Paths => (0 => (I0_ipd'last_event, tpd_I0_O, TRUE),
                 1 => (I1_ipd'last_event, tpd_I1_O, TRUE),
                 2 => (I2_ipd'last_event, tpd_I2_O, TRUE),
                 3 => (I3_ipd'last_event, tpd_I3_O, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;

configuration CFG_NAN4_VITAL of NAN4 is 
        for VITAL_VF
        end for; 
end CFG_NAN4_VITAL;
----- VITAL model for cell NAN5 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity NAN5 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_I0_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I1_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I2_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I3_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I4_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tipd_I0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I2                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I3                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I4                        :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      I0                             :	in    STD_ULOGIC;
      I1                             :	in    STD_ULOGIC;
      I2                             :	in    STD_ULOGIC;
      I3                             :	in    STD_ULOGIC;
      I4                             :	in    STD_ULOGIC;
      O                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of NAN5 : entity is TRUE;
end NAN5;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library VF1;
architecture VITAL_VF of NAN5 is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL I0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I1_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I2_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I3_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I4_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (I0_ipd, I0, tipd_I0);
   VitalWireDelay (I1_ipd, I1, tipd_I1);
   VitalWireDelay (I2_ipd, I2, tipd_I2);
   VitalWireDelay (I3_ipd, I3, tipd_I3);
   VitalWireDelay (I4_ipd, I4, tipd_I4);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (I0_ipd, I1_ipd, I2_ipd, I3_ipd, I4_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS O_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE O_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      O_zd :=
       ((NOT I1_ipd)) OR ((NOT I0_ipd)) OR ((NOT I2_ipd)) OR ((NOT I3_ipd))
         OR ((NOT I4_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => O,
       GlitchData => O_GlitchData,
       OutSignalName => "O",
       OutTemp => O_zd,
       Paths => (0 => (I0_ipd'last_event, tpd_I0_O, TRUE),
                 1 => (I1_ipd'last_event, tpd_I1_O, TRUE),
                 2 => (I2_ipd'last_event, tpd_I2_O, TRUE),
                 3 => (I3_ipd'last_event, tpd_I3_O, TRUE),
                 4 => (I4_ipd'last_event, tpd_I4_O, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;

configuration CFG_NAN5_VITAL of NAN5 is 
        for VITAL_VF
        end for; 
end CFG_NAN5_VITAL;
----- VITAL model for cell NAN6 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity NAN6 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_I0_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I1_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I2_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I3_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I4_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I5_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tipd_I0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I2                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I3                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I4                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I5                        :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      I0                             :	in    STD_ULOGIC;
      I1                             :	in    STD_ULOGIC;
      I2                             :	in    STD_ULOGIC;
      I3                             :	in    STD_ULOGIC;
      I4                             :	in    STD_ULOGIC;
      I5                             :	in    STD_ULOGIC;
      O                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of NAN6 : entity is TRUE;
end NAN6;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
 
library VF1;
architecture VITAL_VF of NAN6 is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL I0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I1_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I2_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I3_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I4_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I5_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (I0_ipd, I0, tipd_I0);
   VitalWireDelay (I1_ipd, I1, tipd_I1);
   VitalWireDelay (I2_ipd, I2, tipd_I2);
   VitalWireDelay (I3_ipd, I3, tipd_I3);
   VitalWireDelay (I4_ipd, I4, tipd_I4);
   VitalWireDelay (I5_ipd, I5, tipd_I5);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (I0_ipd, I1_ipd, I2_ipd, I3_ipd, I4_ipd, I5_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS O_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE O_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      O_zd :=
       ((NOT I1_ipd)) OR ((NOT I0_ipd)) OR ((NOT I2_ipd)) OR ((NOT I3_ipd))
         OR ((NOT I4_ipd)) OR ((NOT I5_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => O,
       GlitchData => O_GlitchData,
       OutSignalName => "O",
       OutTemp => O_zd,
       Paths => (0 => (I0_ipd'last_event, tpd_I0_O, TRUE),
                 1 => (I1_ipd'last_event, tpd_I1_O, TRUE),
                 2 => (I2_ipd'last_event, tpd_I2_O, TRUE),
                 3 => (I3_ipd'last_event, tpd_I3_O, TRUE),
                 4 => (I4_ipd'last_event, tpd_I4_O, TRUE),
                 5 => (I5_ipd'last_event, tpd_I5_O, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;
 
configuration CFG_NAN6_VITAL of NAN6 is 
        for VITAL_VF
        end for; 
end CFG_NAN6_VITAL;
----- VITAL model for cell NAN7 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity NAN7 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_I0_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I1_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I2_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I3_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I4_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I5_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I6_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tipd_I0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I2                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I3                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I4                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I5                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I6                        :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      I0                             :	in    STD_ULOGIC;
      I1                             :	in    STD_ULOGIC;
      I2                             :	in    STD_ULOGIC;
      I3                             :	in    STD_ULOGIC;
      I4                             :	in    STD_ULOGIC;
      I5                             :	in    STD_ULOGIC;
      I6                             :	in    STD_ULOGIC;
      O                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of NAN7 : entity is TRUE;
end NAN7;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
 
library VF1;
architecture VITAL_VF of NAN7 is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL I0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I1_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I2_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I3_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I4_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I5_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I6_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (I0_ipd, I0, tipd_I0);
   VitalWireDelay (I1_ipd, I1, tipd_I1);
   VitalWireDelay (I2_ipd, I2, tipd_I2);
   VitalWireDelay (I3_ipd, I3, tipd_I3);
   VitalWireDelay (I4_ipd, I4, tipd_I4);
   VitalWireDelay (I5_ipd, I5, tipd_I5);
   VitalWireDelay (I6_ipd, I6, tipd_I6);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (I0_ipd, I1_ipd, I2_ipd, I3_ipd, I4_ipd, I5_ipd, I6_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS O_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE O_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      O_zd :=
       ((NOT I1_ipd)) OR ((NOT I0_ipd)) OR ((NOT I2_ipd)) OR ((NOT I3_ipd))
         OR ((NOT I4_ipd)) OR ((NOT I5_ipd)) OR ((NOT I6_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => O,
       GlitchData => O_GlitchData,
       OutSignalName => "O",
       OutTemp => O_zd,
       Paths => (0 => (I0_ipd'last_event, tpd_I0_O, TRUE),
                 1 => (I1_ipd'last_event, tpd_I1_O, TRUE),
                 2 => (I2_ipd'last_event, tpd_I2_O, TRUE),
                 3 => (I3_ipd'last_event, tpd_I3_O, TRUE),
                 4 => (I4_ipd'last_event, tpd_I4_O, TRUE),
                 5 => (I5_ipd'last_event, tpd_I5_O, TRUE),
                 6 => (I6_ipd'last_event, tpd_I6_O, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;
 
configuration CFG_NAN7_VITAL of NAN7 is 
        for VITAL_VF
        end for; 
end CFG_NAN7_VITAL;
----- VITAL model for cell NAN8 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity NAN8 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_I0_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I1_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I2_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I3_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I4_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I5_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I6_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I7_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tipd_I0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I2                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I3                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I4                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I5                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I6                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I7                        :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      I0                             :	in    STD_ULOGIC;
      I1                             :	in    STD_ULOGIC;
      I2                             :	in    STD_ULOGIC;
      I3                             :	in    STD_ULOGIC;
      I4                             :	in    STD_ULOGIC;
      I5                             :	in    STD_ULOGIC;
      I6                             :	in    STD_ULOGIC;
      I7                             :	in    STD_ULOGIC;
      O                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of NAN8 : entity is TRUE;
end NAN8;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
 
library VF1;
architecture VITAL_VF of NAN8 is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL I0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I1_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I2_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I3_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I4_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I5_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I6_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I7_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (I0_ipd, I0, tipd_I0);
   VitalWireDelay (I1_ipd, I1, tipd_I1);
   VitalWireDelay (I2_ipd, I2, tipd_I2);
   VitalWireDelay (I3_ipd, I3, tipd_I3);
   VitalWireDelay (I4_ipd, I4, tipd_I4);
   VitalWireDelay (I5_ipd, I5, tipd_I5);
   VitalWireDelay (I6_ipd, I6, tipd_I6);
   VitalWireDelay (I7_ipd, I7, tipd_I7);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (I0_ipd, I1_ipd, I2_ipd, I3_ipd, I4_ipd, I5_ipd, I6_ipd, I7_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS O_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE O_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      O_zd :=
       ((NOT I1_ipd)) OR ((NOT I0_ipd)) OR ((NOT I2_ipd)) OR ((NOT I3_ipd))
         OR ((NOT I4_ipd)) OR ((NOT I5_ipd)) OR ((NOT I6_ipd)) OR ((NOT
         I7_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => O,
       GlitchData => O_GlitchData,
       OutSignalName => "O",
       OutTemp => O_zd,
       Paths => (0 => (I0_ipd'last_event, tpd_I0_O, TRUE),
                 1 => (I1_ipd'last_event, tpd_I1_O, TRUE),
                 2 => (I2_ipd'last_event, tpd_I2_O, TRUE),
                 3 => (I3_ipd'last_event, tpd_I3_O, TRUE),
                 4 => (I4_ipd'last_event, tpd_I4_O, TRUE),
                 5 => (I5_ipd'last_event, tpd_I5_O, TRUE),
                 6 => (I6_ipd'last_event, tpd_I6_O, TRUE),
                 7 => (I7_ipd'last_event, tpd_I7_O, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;
 
configuration CFG_NAN8_VITAL of NAN8 is 
        for VITAL_VF
        end for; 
end CFG_NAN8_VITAL;
----- VITAL model for cell NEQ22 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity NEQ22 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_A0_O                       :	VitalDelayType01 := (1.800 ns, 1.800 ns);
      tpd_A1_O                       :	VitalDelayType01 := (1.800 ns, 1.800 ns);
      tpd_B0_O                       :	VitalDelayType01 := (1.800 ns, 1.800 ns);
      tpd_B1_O                       :	VitalDelayType01 := (1.800 ns, 1.800 ns);
      tipd_A0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_A1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A0                             :	in    STD_ULOGIC;
      A1                             :	in    STD_ULOGIC;
      B0                             :	in    STD_ULOGIC;
      B1                             :	in    STD_ULOGIC;
      O                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of NEQ22 : entity is TRUE;
end NEQ22;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_VF of NEQ22 is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL A0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL A1_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B1_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A0_ipd, A0, tipd_A0);
   VitalWireDelay (A1_ipd, A1, tipd_A1);
   VitalWireDelay (B0_ipd, B0, tipd_B0);
   VitalWireDelay (B1_ipd, B1, tipd_B1);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A0_ipd, A1_ipd, B0_ipd, B1_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS O_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE O_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      O_zd := ((B1_ipd) XOR (A1_ipd)) OR ((B0_ipd) XOR (A0_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => O,
       GlitchData => O_GlitchData,
       OutSignalName => "O",
       OutTemp => O_zd,
       Paths => (0 => (A0_ipd'last_event, tpd_A0_O, TRUE),
                 1 => (A1_ipd'last_event, tpd_A1_O, TRUE),
                 2 => (B0_ipd'last_event, tpd_B0_O, TRUE),
                 3 => (B1_ipd'last_event, tpd_B1_O, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;

configuration CFG_NEQ22_VITAL of NEQ22 is 
        for VITAL_VF
        end for; 
end CFG_NEQ22_VITAL;
----- VITAL model for cell NOR2 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity NOR2 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_I0_O                       :	VitalDelayType01 := (1.25 ns, 1.25 ns);
      tpd_I1_O                       :	VitalDelayType01 := (1.25 ns, 1.25 ns);
      tipd_I0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      I0                             :	in    STD_ULOGIC;
      I1                             :	in    STD_ULOGIC;
      O                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of NOR2 : entity is TRUE;
end NOR2;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library VF1;
architecture VITAL_VF of NOR2 is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL I0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I1_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (I0_ipd, I0, tipd_I0);
   VitalWireDelay (I1_ipd, I1, tipd_I1);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (I0_ipd, I1_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS O_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE O_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      O_zd := ((NOT I1_ipd)) AND ((NOT I0_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => O,
       GlitchData => O_GlitchData,
       OutSignalName => "O",
       OutTemp => O_zd,
       Paths => (0 => (I0_ipd'last_event, tpd_I0_O, TRUE),
                 1 => (I1_ipd'last_event, tpd_I1_O, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;

configuration CFG_NOR2_VITAL of NOR2 is 
        for VITAL_VF
        end for; 
end CFG_NOR2_VITAL;
----- VITAL model for cell NOR3 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity NOR3 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_I0_O                       :	VitalDelayType01 := (1.25 ns, 1.25 ns);
      tpd_I1_O                       :	VitalDelayType01 := (1.25 ns, 1.25 ns);
      tpd_I2_O                       :	VitalDelayType01 := (1.25 ns, 1.25 ns);
      tipd_I0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I2                        :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      I0                             :	in    STD_ULOGIC;
      I1                             :	in    STD_ULOGIC;
      I2                             :	in    STD_ULOGIC;
      O                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of NOR3 : entity is TRUE;
end NOR3;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library VF1;
architecture VITAL_VF of NOR3 is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL I0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I1_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I2_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (I0_ipd, I0, tipd_I0);
   VitalWireDelay (I1_ipd, I1, tipd_I1);
   VitalWireDelay (I2_ipd, I2, tipd_I2);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (I0_ipd, I1_ipd, I2_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS O_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE O_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      O_zd := ((NOT I1_ipd)) AND ((NOT I0_ipd)) AND ((NOT I2_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => O,
       GlitchData => O_GlitchData,
       OutSignalName => "O",
       OutTemp => O_zd,
       Paths => (0 => (I0_ipd'last_event, tpd_I0_O, TRUE),
                 1 => (I1_ipd'last_event, tpd_I1_O, TRUE),
                 2 => (I2_ipd'last_event, tpd_I2_O, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;

configuration CFG_NOR3_VITAL of NOR3 is 
        for VITAL_VF
        end for; 
end CFG_NOR3_VITAL;
----- VITAL model for cell NOR4 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity NOR4 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_I0_O                       :	VitalDelayType01 := (1.80 ns, 1.80 ns);
      tpd_I1_O                       :	VitalDelayType01 := (1.80 ns, 1.80 ns);
      tpd_I2_O                       :	VitalDelayType01 := (1.80 ns, 1.80 ns);
      tpd_I3_O                       :	VitalDelayType01 := (1.80 ns, 1.80 ns);
      tipd_I0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I2                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I3                        :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      I0                             :	in    STD_ULOGIC;
      I1                             :	in    STD_ULOGIC;
      I2                             :	in    STD_ULOGIC;
      I3                             :	in    STD_ULOGIC;
      O                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of NOR4 : entity is TRUE;
end NOR4;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library VF1;
architecture VITAL_VF of NOR4 is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL I0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I1_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I2_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I3_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (I0_ipd, I0, tipd_I0);
   VitalWireDelay (I1_ipd, I1, tipd_I1);
   VitalWireDelay (I2_ipd, I2, tipd_I2);
   VitalWireDelay (I3_ipd, I3, tipd_I3);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (I0_ipd, I1_ipd, I2_ipd, I3_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS O_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE O_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      O_zd :=
       ((NOT I1_ipd)) AND ((NOT I0_ipd)) AND ((NOT I2_ipd)) AND ((NOT
         I3_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => O,
       GlitchData => O_GlitchData,
       OutSignalName => "O",
       OutTemp => O_zd,
       Paths => (0 => (I0_ipd'last_event, tpd_I0_O, TRUE),
                 1 => (I1_ipd'last_event, tpd_I1_O, TRUE),
                 2 => (I2_ipd'last_event, tpd_I2_O, TRUE),
                 3 => (I3_ipd'last_event, tpd_I3_O, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;

configuration CFG_NOR4_VITAL of NOR4 is 
        for VITAL_VF
        end for; 
end CFG_NOR4_VITAL;
----- VITAL model for cell NOR5 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity NOR5 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_I0_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I1_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I2_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I3_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I4_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tipd_I0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I2                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I3                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I4                        :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      I0                             :	in    STD_ULOGIC;
      I1                             :	in    STD_ULOGIC;
      I2                             :	in    STD_ULOGIC;
      I3                             :	in    STD_ULOGIC;
      I4                             :	in    STD_ULOGIC;
      O                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of NOR5 : entity is TRUE;
end NOR5;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
 
library VF1;
architecture VITAL_VF of NOR5 is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL I0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I1_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I2_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I3_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I4_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (I0_ipd, I0, tipd_I0);
   VitalWireDelay (I1_ipd, I1, tipd_I1);
   VitalWireDelay (I2_ipd, I2, tipd_I2);
   VitalWireDelay (I3_ipd, I3, tipd_I3);
   VitalWireDelay (I4_ipd, I4, tipd_I4);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (I0_ipd, I1_ipd, I2_ipd, I3_ipd, I4_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS O_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE O_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      O_zd :=
       ((NOT I1_ipd)) AND ((NOT I0_ipd)) AND ((NOT I2_ipd)) AND ((NOT
         I3_ipd)) AND ((NOT I4_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => O,
       GlitchData => O_GlitchData,
       OutSignalName => "O",
       OutTemp => O_zd,
       Paths => (0 => (I0_ipd'last_event, tpd_I0_O, TRUE),
                 1 => (I1_ipd'last_event, tpd_I1_O, TRUE),
                 2 => (I2_ipd'last_event, tpd_I2_O, TRUE),
                 3 => (I3_ipd'last_event, tpd_I3_O, TRUE),
                 4 => (I4_ipd'last_event, tpd_I4_O, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;
 
configuration CFG_NOR5_VITAL of NOR5 is 
        for VITAL_VF
        end for; 
end CFG_NOR5_VITAL;
----- VITAL model for cell NOR6 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity NOR6 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_I0_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I1_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I2_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I3_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I4_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I5_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tipd_I0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I2                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I3                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I4                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I5                        :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      I0                             :	in    STD_ULOGIC;
      I1                             :	in    STD_ULOGIC;
      I2                             :	in    STD_ULOGIC;
      I3                             :	in    STD_ULOGIC;
      I4                             :	in    STD_ULOGIC;
      I5                             :	in    STD_ULOGIC;
      O                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of NOR6 : entity is TRUE;
end NOR6;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
 
library VF1;
architecture VITAL_VF of NOR6 is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL I0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I1_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I2_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I3_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I4_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I5_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (I0_ipd, I0, tipd_I0);
   VitalWireDelay (I1_ipd, I1, tipd_I1);
   VitalWireDelay (I2_ipd, I2, tipd_I2);
   VitalWireDelay (I3_ipd, I3, tipd_I3);
   VitalWireDelay (I4_ipd, I4, tipd_I4);
   VitalWireDelay (I5_ipd, I5, tipd_I5);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (I0_ipd, I1_ipd, I2_ipd, I3_ipd, I4_ipd, I5_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS O_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE O_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      O_zd :=
       ((NOT I1_ipd)) AND ((NOT I0_ipd)) AND ((NOT I2_ipd)) AND ((NOT
         I3_ipd)) AND ((NOT I4_ipd)) AND ((NOT I5_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => O,
       GlitchData => O_GlitchData,
       OutSignalName => "O",
       OutTemp => O_zd,
       Paths => (0 => (I0_ipd'last_event, tpd_I0_O, TRUE),
                 1 => (I1_ipd'last_event, tpd_I1_O, TRUE),
                 2 => (I2_ipd'last_event, tpd_I2_O, TRUE),
                 3 => (I3_ipd'last_event, tpd_I3_O, TRUE),
                 4 => (I4_ipd'last_event, tpd_I4_O, TRUE),
                 5 => (I5_ipd'last_event, tpd_I5_O, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;
 
configuration CFG_NOR6_VITAL of NOR6 is 
        for VITAL_VF
        end for; 
end CFG_NOR6_VITAL;
----- VITAL model for cell NOR7 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity NOR7 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_I0_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I1_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I2_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I3_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I4_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I5_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I6_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tipd_I0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I2                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I3                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I4                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I5                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I6                        :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      I0                             :	in    STD_ULOGIC;
      I1                             :	in    STD_ULOGIC;
      I2                             :	in    STD_ULOGIC;
      I3                             :	in    STD_ULOGIC;
      I4                             :	in    STD_ULOGIC;
      I5                             :	in    STD_ULOGIC;
      I6                             :	in    STD_ULOGIC;
      O                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of NOR7 : entity is TRUE;
end NOR7;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
 
library VF1;
architecture VITAL_VF of NOR7 is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL I0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I1_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I2_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I3_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I4_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I5_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I6_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (I0_ipd, I0, tipd_I0);
   VitalWireDelay (I1_ipd, I1, tipd_I1);
   VitalWireDelay (I2_ipd, I2, tipd_I2);
   VitalWireDelay (I3_ipd, I3, tipd_I3);
   VitalWireDelay (I4_ipd, I4, tipd_I4);
   VitalWireDelay (I5_ipd, I5, tipd_I5);
   VitalWireDelay (I6_ipd, I6, tipd_I6);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (I0_ipd, I1_ipd, I2_ipd, I3_ipd, I4_ipd, I5_ipd, I6_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS O_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE O_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      O_zd :=
       ((NOT I1_ipd)) AND ((NOT I0_ipd)) AND ((NOT I2_ipd)) AND ((NOT
         I3_ipd)) AND ((NOT I4_ipd)) AND ((NOT I5_ipd)) AND ((NOT I6_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => O,
       GlitchData => O_GlitchData,
       OutSignalName => "O",
       OutTemp => O_zd,
       Paths => (0 => (I0_ipd'last_event, tpd_I0_O, TRUE),
                 1 => (I1_ipd'last_event, tpd_I1_O, TRUE),
                 2 => (I2_ipd'last_event, tpd_I2_O, TRUE),
                 3 => (I3_ipd'last_event, tpd_I3_O, TRUE),
                 4 => (I4_ipd'last_event, tpd_I4_O, TRUE),
                 5 => (I5_ipd'last_event, tpd_I5_O, TRUE),
                 6 => (I6_ipd'last_event, tpd_I6_O, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;
 
configuration CFG_NOR7_VITAL of NOR7 is 
        for VITAL_VF
        end for; 
end CFG_NOR7_VITAL;
----- VITAL model for cell NOR8 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity NOR8 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_I0_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I1_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I2_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I3_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I4_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I5_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I6_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I7_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tipd_I0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I2                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I3                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I4                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I5                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I6                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I7                        :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      I0                             :	in    STD_ULOGIC;
      I1                             :	in    STD_ULOGIC;
      I2                             :	in    STD_ULOGIC;
      I3                             :	in    STD_ULOGIC;
      I4                             :	in    STD_ULOGIC;
      I5                             :	in    STD_ULOGIC;
      I6                             :	in    STD_ULOGIC;
      I7                             :	in    STD_ULOGIC;
      O                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of NOR8 : entity is TRUE;
end NOR8;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
 
library VF1;
architecture VITAL_VF of NOR8 is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL I0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I1_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I2_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I3_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I4_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I5_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I6_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I7_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (I0_ipd, I0, tipd_I0);
   VitalWireDelay (I1_ipd, I1, tipd_I1);
   VitalWireDelay (I2_ipd, I2, tipd_I2);
   VitalWireDelay (I3_ipd, I3, tipd_I3);
   VitalWireDelay (I4_ipd, I4, tipd_I4);
   VitalWireDelay (I5_ipd, I5, tipd_I5);
   VitalWireDelay (I6_ipd, I6, tipd_I6);
   VitalWireDelay (I7_ipd, I7, tipd_I7);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (I0_ipd, I1_ipd, I2_ipd, I3_ipd, I4_ipd, I5_ipd, I6_ipd, I7_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS O_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE O_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      O_zd :=
       ((NOT I1_ipd)) AND ((NOT I0_ipd)) AND ((NOT I2_ipd)) AND ((NOT
         I3_ipd)) AND ((NOT I4_ipd)) AND ((NOT I5_ipd)) AND ((NOT I6_ipd))
         AND ((NOT I7_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => O,
       GlitchData => O_GlitchData,
       OutSignalName => "O",
       OutTemp => O_zd,
       Paths => (0 => (I0_ipd'last_event, tpd_I0_O, TRUE),
                 1 => (I1_ipd'last_event, tpd_I1_O, TRUE),
                 2 => (I2_ipd'last_event, tpd_I2_O, TRUE),
                 3 => (I3_ipd'last_event, tpd_I3_O, TRUE),
                 4 => (I4_ipd'last_event, tpd_I4_O, TRUE),
                 5 => (I5_ipd'last_event, tpd_I5_O, TRUE),
                 6 => (I6_ipd'last_event, tpd_I6_O, TRUE),
                 7 => (I7_ipd'last_event, tpd_I7_O, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;
 
configuration CFG_NOR8_VITAL of NOR8 is 
        for VITAL_VF
        end for; 
end CFG_NOR8_VITAL;
----- VITAL model for cell OA21 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity OA21 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_I0_O                       :	VitalDelayType01 := (1.25 ns, 1.25 ns);
      tpd_I1_O                       :	VitalDelayType01 := (1.25 ns, 1.25 ns);
      tpd_I2_O                       :	VitalDelayType01 := (1.25 ns, 1.25 ns);
      tipd_I0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I2                        :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      I0                             :	in    STD_ULOGIC;
      I1                             :	in    STD_ULOGIC;
      I2                             :	in    STD_ULOGIC;
      O                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of OA21 : entity is TRUE;
end OA21;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library VF1;
architecture VITAL_VF of OA21 is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL I0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I1_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I2_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (I0_ipd, I0, tipd_I0);
   VitalWireDelay (I1_ipd, I1, tipd_I1);
   VitalWireDelay (I2_ipd, I2, tipd_I2);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (I0_ipd, I1_ipd, I2_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS O_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE O_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      O_zd := (I2_ipd) AND ((I1_ipd) OR (I0_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => O,
       GlitchData => O_GlitchData,
       OutSignalName => "O",
       OutTemp => O_zd,
       Paths => (0 => (I0_ipd'last_event, tpd_I0_O, TRUE),
                 1 => (I1_ipd'last_event, tpd_I1_O, TRUE),
                 2 => (I2_ipd'last_event, tpd_I2_O, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;

configuration CFG_OA21_VITAL of OA21 is 
        for VITAL_VF
        end for; 
end CFG_OA21_VITAL;
----- VITAL model for cell OA221 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity OA221 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_I0_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I1_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I2_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I3_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I4_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tipd_I0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I2                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I3                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I4                        :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      I0                             :	in    STD_ULOGIC;
      I1                             :	in    STD_ULOGIC;
      I2                             :	in    STD_ULOGIC;
      I3                             :	in    STD_ULOGIC;
      I4                             :	in    STD_ULOGIC;
      O                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of OA221 : entity is TRUE;
end OA221;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
 
library VF1;
architecture VITAL_VF of OA221 is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL I0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I1_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I2_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I3_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I4_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (I0_ipd, I0, tipd_I0);
   VitalWireDelay (I1_ipd, I1, tipd_I1);
   VitalWireDelay (I2_ipd, I2, tipd_I2);
   VitalWireDelay (I3_ipd, I3, tipd_I3);
   VitalWireDelay (I4_ipd, I4, tipd_I4);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (I0_ipd, I1_ipd, I2_ipd, I3_ipd, I4_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS O_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE O_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      O_zd :=
       ((I3_ipd) OR (I2_ipd)) AND ((I1_ipd) OR (I0_ipd)) AND (I4_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => O,
       GlitchData => O_GlitchData,
       OutSignalName => "O",
       OutTemp => O_zd,
       Paths => (0 => (I0_ipd'last_event, tpd_I0_O, TRUE),
                 1 => (I1_ipd'last_event, tpd_I1_O, TRUE),
                 2 => (I2_ipd'last_event, tpd_I2_O, TRUE),
                 3 => (I3_ipd'last_event, tpd_I3_O, TRUE),
                 4 => (I4_ipd'last_event, tpd_I4_O, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;
 
configuration CFG_OA221_VITAL of OA221 is 
        for VITAL_VF
        end for; 
end CFG_OA221_VITAL;
----- VITAL model for cell OA321 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity OA321 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_I0_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I1_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I2_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I3_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I4_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I5_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tipd_I0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I2                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I3                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I4                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I5                        :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      I0                             :	in    STD_ULOGIC;
      I1                             :	in    STD_ULOGIC;
      I2                             :	in    STD_ULOGIC;
      I3                             :	in    STD_ULOGIC;
      I4                             :	in    STD_ULOGIC;
      I5                             :	in    STD_ULOGIC;
      O                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of OA321 : entity is TRUE;
end OA321;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
 
library VF1;
architecture VITAL_VF of OA321 is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL I0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I1_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I2_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I3_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I4_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I5_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (I0_ipd, I0, tipd_I0);
   VitalWireDelay (I1_ipd, I1, tipd_I1);
   VitalWireDelay (I2_ipd, I2, tipd_I2);
   VitalWireDelay (I3_ipd, I3, tipd_I3);
   VitalWireDelay (I4_ipd, I4, tipd_I4);
   VitalWireDelay (I5_ipd, I5, tipd_I5);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (I0_ipd, I1_ipd, I2_ipd, I3_ipd, I4_ipd, I5_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS O_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE O_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      O_zd :=
       ((I4_ipd) OR (I3_ipd)) AND ((I1_ipd) OR (I0_ipd) OR (I2_ipd)) AND
         (I5_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => O,
       GlitchData => O_GlitchData,
       OutSignalName => "O",
       OutTemp => O_zd,
       Paths => (0 => (I0_ipd'last_event, tpd_I0_O, TRUE),
                 1 => (I1_ipd'last_event, tpd_I1_O, TRUE),
                 2 => (I2_ipd'last_event, tpd_I2_O, TRUE),
                 3 => (I3_ipd'last_event, tpd_I3_O, TRUE),
                 4 => (I4_ipd'last_event, tpd_I4_O, TRUE),
                 5 => (I5_ipd'last_event, tpd_I5_O, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;
 
configuration CFG_OA321_VITAL of OA321 is 
        for VITAL_VF
        end for; 
end CFG_OA321_VITAL;
----- VITAL model for cell OBUF -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;

LIBRARY VF1 ;
use VF1.VLOGTOVITAL_TABLES.all;



-- entity declaration --
entity OBUF is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_I0_O                       :	VitalDelayType01 := (1.70 ns, 1.70 ns);
      tipd_I0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      I0                             :	in    STD_ULOGIC;
      O                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of OBUF : entity is TRUE;
end OBUF;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library VF1;
-- use VF1.VTABLES.all;
architecture VITAL_VF of OBUF is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL I0_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (I0_ipd, I0, tipd_I0);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (I0_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS O_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE O_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      O_zd := TO_X01(I0_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => O,
       GlitchData => O_GlitchData,
       OutSignalName => "O",
       OutTemp => O_zd,
       Paths => (0 => (I0_ipd'last_event, tpd_I0_O, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;

configuration CFG_OBUF_VITAL of OBUF is 
        for VITAL_VF
        end for; 
end CFG_OBUF_VITAL;

----- VITAL model for cell OR2 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity OR2 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_I0_O                       :	VitalDelayType01 := (1.25 ns, 1.25 ns);
      tpd_I1_O                       :	VitalDelayType01 := (1.25 ns, 1.25 ns);
      tipd_I0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      I0                             :	in    STD_ULOGIC;
      I1                             :	in    STD_ULOGIC;
      O                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of OR2 : entity is TRUE;
end OR2;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library VF1;
architecture VITAL_VF of OR2 is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL I0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I1_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (I0_ipd, I0, tipd_I0);
   VitalWireDelay (I1_ipd, I1, tipd_I1);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (I0_ipd, I1_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS O_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE O_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      O_zd := (I1_ipd) OR (I0_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => O,
       GlitchData => O_GlitchData,
       OutSignalName => "O",
       OutTemp => O_zd,
       Paths => (0 => (I0_ipd'last_event, tpd_I0_O, TRUE),
                 1 => (I1_ipd'last_event, tpd_I1_O, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;

configuration CFG_OR2_VITAL of OR2 is 
        for VITAL_VF
        end for; 
end CFG_OR2_VITAL;
----- VITAL model for cell OR3 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity OR3 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_I0_O                       :	VitalDelayType01 := (1.25 ns, 1.25 ns);
      tpd_I1_O                       :	VitalDelayType01 := (1.25 ns, 1.25 ns);
      tpd_I2_O                       :	VitalDelayType01 := (1.25 ns, 1.25 ns);
      tipd_I0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I2                        :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      I0                             :	in    STD_ULOGIC;
      I1                             :	in    STD_ULOGIC;
      I2                             :	in    STD_ULOGIC;
      O                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of OR3 : entity is TRUE;
end OR3;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library VF1;
architecture VITAL_VF of OR3 is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL I0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I1_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I2_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (I0_ipd, I0, tipd_I0);
   VitalWireDelay (I1_ipd, I1, tipd_I1);
   VitalWireDelay (I2_ipd, I2, tipd_I2);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (I0_ipd, I1_ipd, I2_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS O_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE O_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      O_zd := (I1_ipd) OR (I0_ipd) OR (I2_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => O,
       GlitchData => O_GlitchData,
       OutSignalName => "O",
       OutTemp => O_zd,
       Paths => (0 => (I0_ipd'last_event, tpd_I0_O, TRUE),
                 1 => (I1_ipd'last_event, tpd_I1_O, TRUE),
                 2 => (I2_ipd'last_event, tpd_I2_O, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;

configuration CFG_OR3_VITAL of OR3 is 
        for VITAL_VF
        end for; 
end CFG_OR3_VITAL;
----- VITAL model for cell OR4 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity OR4 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_I0_O                       :	VitalDelayType01 := (1.80 ns, 1.80 ns);
      tpd_I1_O                       :	VitalDelayType01 := (1.80 ns, 1.80 ns);
      tpd_I2_O                       :	VitalDelayType01 := (1.80 ns, 1.80 ns);
      tpd_I3_O                       :	VitalDelayType01 := (1.80 ns, 1.80 ns);
      tipd_I0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I2                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I3                        :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      I0                             :	in    STD_ULOGIC;
      I1                             :	in    STD_ULOGIC;
      I2                             :	in    STD_ULOGIC;
      I3                             :	in    STD_ULOGIC;
      O                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of OR4 : entity is TRUE;
end OR4;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library VF1;
architecture VITAL_VF of OR4 is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL I0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I1_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I2_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I3_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (I0_ipd, I0, tipd_I0);
   VitalWireDelay (I1_ipd, I1, tipd_I1);
   VitalWireDelay (I2_ipd, I2, tipd_I2);
   VitalWireDelay (I3_ipd, I3, tipd_I3);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (I0_ipd, I1_ipd, I2_ipd, I3_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS O_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE O_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      O_zd := (I1_ipd) OR (I0_ipd) OR (I2_ipd) OR (I3_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => O,
       GlitchData => O_GlitchData,
       OutSignalName => "O",
       OutTemp => O_zd,
       Paths => (0 => (I0_ipd'last_event, tpd_I0_O, TRUE),
                 1 => (I1_ipd'last_event, tpd_I1_O, TRUE),
                 2 => (I2_ipd'last_event, tpd_I2_O, TRUE),
                 3 => (I3_ipd'last_event, tpd_I3_O, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;

configuration CFG_OR4_VITAL of OR4 is 
        for VITAL_VF
        end for; 
end CFG_OR4_VITAL;
----- VITAL model for cell OR5 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity OR5 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_I0_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I1_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I2_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I3_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I4_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tipd_I0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I2                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I3                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I4                        :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      I0                             :	in    STD_ULOGIC;
      I1                             :	in    STD_ULOGIC;
      I2                             :	in    STD_ULOGIC;
      I3                             :	in    STD_ULOGIC;
      I4                             :	in    STD_ULOGIC;
      O                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of OR5 : entity is TRUE;
end OR5;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
 
library VF1;
architecture VITAL_VF of OR5 is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL I0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I1_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I2_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I3_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I4_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (I0_ipd, I0, tipd_I0);
   VitalWireDelay (I1_ipd, I1, tipd_I1);
   VitalWireDelay (I2_ipd, I2, tipd_I2);
   VitalWireDelay (I3_ipd, I3, tipd_I3);
   VitalWireDelay (I4_ipd, I4, tipd_I4);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (I0_ipd, I1_ipd, I2_ipd, I3_ipd, I4_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS O_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE O_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      O_zd := (I1_ipd) OR (I0_ipd) OR (I2_ipd) OR (I3_ipd) OR (I4_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => O,
       GlitchData => O_GlitchData,
       OutSignalName => "O",
       OutTemp => O_zd,
       Paths => (0 => (I0_ipd'last_event, tpd_I0_O, TRUE),
                 1 => (I1_ipd'last_event, tpd_I1_O, TRUE),
                 2 => (I2_ipd'last_event, tpd_I2_O, TRUE),
                 3 => (I3_ipd'last_event, tpd_I3_O, TRUE),
                 4 => (I4_ipd'last_event, tpd_I4_O, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;
 
configuration CFG_OR5_VITAL of OR5 is 
        for VITAL_VF
        end for; 
end CFG_OR5_VITAL;
----- VITAL model for cell OR6 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity OR6 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_I0_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I1_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I2_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I3_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I4_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I5_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tipd_I0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I2                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I3                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I4                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I5                        :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      I0                             :	in    STD_ULOGIC;
      I1                             :	in    STD_ULOGIC;
      I2                             :	in    STD_ULOGIC;
      I3                             :	in    STD_ULOGIC;
      I4                             :	in    STD_ULOGIC;
      I5                             :	in    STD_ULOGIC;
      O                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of OR6 : entity is TRUE;
end OR6;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
 
library VF1;
architecture VITAL_VF of OR6 is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL I0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I1_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I2_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I3_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I4_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I5_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (I0_ipd, I0, tipd_I0);
   VitalWireDelay (I1_ipd, I1, tipd_I1);
   VitalWireDelay (I2_ipd, I2, tipd_I2);
   VitalWireDelay (I3_ipd, I3, tipd_I3);
   VitalWireDelay (I4_ipd, I4, tipd_I4);
   VitalWireDelay (I5_ipd, I5, tipd_I5);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (I0_ipd, I1_ipd, I2_ipd, I3_ipd, I4_ipd, I5_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS O_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE O_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      O_zd :=
       (I1_ipd) OR (I0_ipd) OR (I2_ipd) OR (I3_ipd) OR (I4_ipd) OR (I5_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => O,
       GlitchData => O_GlitchData,
       OutSignalName => "O",
       OutTemp => O_zd,
       Paths => (0 => (I0_ipd'last_event, tpd_I0_O, TRUE),
                 1 => (I1_ipd'last_event, tpd_I1_O, TRUE),
                 2 => (I2_ipd'last_event, tpd_I2_O, TRUE),
                 3 => (I3_ipd'last_event, tpd_I3_O, TRUE),
                 4 => (I4_ipd'last_event, tpd_I4_O, TRUE),
                 5 => (I5_ipd'last_event, tpd_I5_O, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;
 
configuration CFG_OR6_VITAL of OR6 is 
        for VITAL_VF
        end for; 
end CFG_OR6_VITAL;
----- VITAL model for cell OR7 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity OR7 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_I0_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I1_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I2_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I3_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I4_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I5_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I6_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tipd_I0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I2                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I3                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I4                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I5                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I6                        :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      I0                             :	in    STD_ULOGIC;
      I1                             :	in    STD_ULOGIC;
      I2                             :	in    STD_ULOGIC;
      I3                             :	in    STD_ULOGIC;
      I4                             :	in    STD_ULOGIC;
      I5                             :	in    STD_ULOGIC;
      I6                             :	in    STD_ULOGIC;
      O                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of OR7 : entity is TRUE;
end OR7;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
 
library VF1;
architecture VITAL_VF of OR7 is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL I0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I1_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I2_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I3_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I4_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I5_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I6_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (I0_ipd, I0, tipd_I0);
   VitalWireDelay (I1_ipd, I1, tipd_I1);
   VitalWireDelay (I2_ipd, I2, tipd_I2);
   VitalWireDelay (I3_ipd, I3, tipd_I3);
   VitalWireDelay (I4_ipd, I4, tipd_I4);
   VitalWireDelay (I5_ipd, I5, tipd_I5);
   VitalWireDelay (I6_ipd, I6, tipd_I6);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (I0_ipd, I1_ipd, I2_ipd, I3_ipd, I4_ipd, I5_ipd, I6_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS O_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE O_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      O_zd :=
       (I1_ipd) OR (I0_ipd) OR (I2_ipd) OR (I3_ipd) OR (I4_ipd) OR (I5_ipd)
         OR (I6_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => O,
       GlitchData => O_GlitchData,
       OutSignalName => "O",
       OutTemp => O_zd,
       Paths => (0 => (I0_ipd'last_event, tpd_I0_O, TRUE),
                 1 => (I1_ipd'last_event, tpd_I1_O, TRUE),
                 2 => (I2_ipd'last_event, tpd_I2_O, TRUE),
                 3 => (I3_ipd'last_event, tpd_I3_O, TRUE),
                 4 => (I4_ipd'last_event, tpd_I4_O, TRUE),
                 5 => (I5_ipd'last_event, tpd_I5_O, TRUE),
                 6 => (I6_ipd'last_event, tpd_I6_O, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;
 
configuration CFG_OR7_VITAL of OR7 is 
        for VITAL_VF
        end for; 
end CFG_OR7_VITAL;
----- VITAL model for cell OR8 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity OR8 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_I0_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I1_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I2_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I3_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I4_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I5_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I6_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I7_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tipd_I0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I2                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I3                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I4                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I5                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I6                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I7                        :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      I0                             :	in    STD_ULOGIC;
      I1                             :	in    STD_ULOGIC;
      I2                             :	in    STD_ULOGIC;
      I3                             :	in    STD_ULOGIC;
      I4                             :	in    STD_ULOGIC;
      I5                             :	in    STD_ULOGIC;
      I6                             :	in    STD_ULOGIC;
      I7                             :	in    STD_ULOGIC;
      O                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of OR8 : entity is TRUE;
end OR8;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
 
library VF1;
architecture VITAL_VF of OR8 is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL I0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I1_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I2_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I3_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I4_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I5_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I6_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I7_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (I0_ipd, I0, tipd_I0);
   VitalWireDelay (I1_ipd, I1, tipd_I1);
   VitalWireDelay (I2_ipd, I2, tipd_I2);
   VitalWireDelay (I3_ipd, I3, tipd_I3);
   VitalWireDelay (I4_ipd, I4, tipd_I4);
   VitalWireDelay (I5_ipd, I5, tipd_I5);
   VitalWireDelay (I6_ipd, I6, tipd_I6);
   VitalWireDelay (I7_ipd, I7, tipd_I7);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (I0_ipd, I1_ipd, I2_ipd, I3_ipd, I4_ipd, I5_ipd, I6_ipd, I7_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS O_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE O_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      O_zd :=
       (I1_ipd) OR (I0_ipd) OR (I2_ipd) OR (I3_ipd) OR (I4_ipd) OR (I5_ipd)
         OR (I6_ipd) OR (I7_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => O,
       GlitchData => O_GlitchData,
       OutSignalName => "O",
       OutTemp => O_zd,
       Paths => (0 => (I0_ipd'last_event, tpd_I0_O, TRUE),
                 1 => (I1_ipd'last_event, tpd_I1_O, TRUE),
                 2 => (I2_ipd'last_event, tpd_I2_O, TRUE),
                 3 => (I3_ipd'last_event, tpd_I3_O, TRUE),
                 4 => (I4_ipd'last_event, tpd_I4_O, TRUE),
                 5 => (I5_ipd'last_event, tpd_I5_O, TRUE),
                 6 => (I6_ipd'last_event, tpd_I6_O, TRUE),
                 7 => (I7_ipd'last_event, tpd_I7_O, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;
 
configuration CFG_OR8_VITAL of OR8 is 
        for VITAL_VF
        end for; 
end CFG_OR8_VITAL;
----- VITAL model for cell PUC -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity PUC is
attribute VITAL_LEVEL0 of PUC : entity is TRUE;
end PUC;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library VF1;
architecture VITAL_VF of PUC is
   attribute VITAL_LEVEL0 of VITAL_VF : architecture is TRUE;


begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   --  empty
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------


end VITAL_VF;

configuration CFG_PUC_VITAL of PUC is 
        for VITAL_VF
        end for; 
end CFG_PUC_VITAL;
----- VITAL model for cell RBC -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity RBC is
attribute VITAL_LEVEL0 of RBC : entity is TRUE;
end RBC;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library VF1;
architecture VITAL_VF of RBC is
   attribute VITAL_LEVEL0 of VITAL_VF : architecture is TRUE;


begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   --  empty
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------


end VITAL_VF;

configuration CFG_RBC_VITAL of RBC is 
        for VITAL_VF
        end for; 
end CFG_RBC_VITAL;
----- VITAL model for cell RI -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;

LIBRARY VF1 ;
use VF1.VLOGTOVITAL_TABLES.all;


-- entity declaration --
entity RI is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_CLK_Q                      :	VitalDelayType01 := (1.230 ns, 1.230 ns);
      tsetup_D_CLK_noedge_posedge    :	VitalDelayType := 0.000 ns;---0.330 ns;
      thold_D_CLK_noedge_posedge     :	VitalDelayType := 0.530 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 1.320 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.660 ns;
      ticd_CLK                       :	VitalDelayType := 0.000 ns;
      tisd_D_CLK                     :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of RI : entity is TRUE;
end RI;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library VF1;
architecture VITAL_VF of RI is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL D_CLK_dly	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   VitalSignalDelay (CLK_dly, CLK_ipd, ticd_CLK);
   VitalSignalDelay (D_CLK_dly, D_ipd, tisd_D_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (CLK_dly, D_CLK_dly)

   -- timing check results
   VARIABLE Tviol_D_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 3);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_posedge,
          TimingData              => Tmkr_D_CLK_posedge,
          TestSignal              => D_CLK_dly,
          TestSignalName          => "D",
          TestDelay               => tisd_D_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          SetupHigh               => tsetup_D_CLK_noedge_posedge,
          SetupLow                => tsetup_D_CLK_noedge_posedge,
          HoldHigh                => thold_D_CLK_noedge_posedge,
          HoldLow                 => thold_D_CLK_noedge_posedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/RI",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_dly,
          TestSignalName          => "CLK",
          TestDelay               => ticd_CLK,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/RI",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_posedge or Pviol_CLK;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => dfftab,
        DataIn => (
               D_CLK_dly, CLK_dly, '1','1'));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (CLK_dly'last_event, tpd_CLK_Q, TRUE)),
       Mode => VitalInertial,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;

configuration CFG_RI_VITAL of RI is 
        for VITAL_VF
        end for; 
end CFG_RI_VITAL;
----- VITAL model for cell RIR -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;

LIBRARY VF1 ;
use VF1.VLOGTOVITAL_TABLES.all;



-- entity declaration --
entity RIR is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_R_Q                        :	VitalDelayType01 := (1.230 ns, 1.230 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.230 ns, 1.230 ns);
      tsetup_D_CLK_noedge_posedge :	VitalDelayType := 0.000 ns;---0.330 ns;
      thold_D_CLK_noedge_posedge :	VitalDelayType := 0.530 ns;
      tpw_CLK_posedge         :	VitalDelayType := 0.660 ns;
      tperiod_CLK_posedge             :	VitalDelayType := 1.320 ns;
      trecovery_R_CLK_posedge_posedge :	VitalDelayType := 0.000 ns;---0.330 ns;
      thold_R_CLK_posedge_posedge    :	VitalDelayType := 0.530 ns;
      ticd_CLK                       :	VitalDelayType := 0.000 ns;
      tisd_D_CLK                     :	VitalDelayType := 0.000 ns;
      tisd_R_CLK                     :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_R                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      R                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of RIR : entity is TRUE;
end RIR;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library VF1;
architecture VITAL_VF of RIR is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL R_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL D_CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL R_CLK_dly	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (R_ipd, R, tipd_R);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   VitalSignalDelay (CLK_dly, CLK_ipd, ticd_CLK);
   VitalSignalDelay (D_CLK_dly, D_ipd, tisd_D_CLK);
   VitalSignalDelay (R_CLK_dly, R_ipd, tisd_R_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (CLK_dly, D_CLK_dly, R_CLK_dly)

   -- timing check results
   VARIABLE Tviol_D_CLK_R_EQ_1_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_R_EQ_1_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_R_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_R_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK_R_EQ_1	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK_R_EQ_1	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 3);
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_R_EQ_1_posedge,
          TimingData              => Tmkr_D_CLK_R_EQ_1_posedge,
          TestSignal              => D_CLK_dly,
          TestSignalName          => "D",
          TestDelay               => tisd_D_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          SetupHigh               => tsetup_D_CLK_noedge_posedge,
          SetupLow                => tsetup_D_CLK_noedge_posedge,
          HoldHigh                => thold_D_CLK_noedge_posedge,
          HoldLow                 => thold_D_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(R_CLK_dly) = '0',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/RIR",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);

         VitalRecoveryRemovalCheck (
          Violation               => Tviol_R_CLK_posedge,
          TimingData              => Tmkr_R_CLK_posedge,
          TestSignal              => R_CLK_dly,
          TestSignalName          => "R",
          TestDelay               => tisd_R_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          Recovery                => trecovery_R_CLK_posedge_posedge,
          Removal                 => thold_R_CLK_posedge_posedge,
          ActiveLow               => FALSE,
          CheckEnabled            => TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/RIR",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK_R_EQ_1,
          PeriodData              => PInfo_CLK_R_EQ_1,
          TestSignal              => CLK_dly,
          TestSignalName          => "CLK",
          TestDelay               => ticd_CLK,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TO_X01((R_CLK_dly) ) = '0',
          HeaderMsg               => InstancePath & "/RIR",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_R_EQ_1_posedge or Tviol_R_CLK_posedge or Pviol_CLK_R_EQ_1;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => dfftab,
        DataIn => (
               D_CLK_dly, CLK_dly,NOT(R_CLK_dly), '1'));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (R_CLK_dly'last_event, tpd_R_Q, TRUE),
                 1 => (CLK_dly'last_event, tpd_CLK_Q, TRUE)),
       Mode => VitalInertial,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;

configuration CFG_RIR_VITAL of RIR is 
        for VITAL_VF
        end for; 
end CFG_RIR_VITAL;
----- VITAL model for cell RIS -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;

LIBRARY VF1 ;
use VF1.VLOGTOVITAL_TABLES.all;



-- entity declaration --
entity RIS is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_S_Q                        :	VitalDelayType01 := (1.230 ns, 1.230 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.230 ns, 1.230 ns);
      tsetup_D_CLK_noedge_posedge :	VitalDelayType := 0.000 ns;---0.330 ns;
      thold_D_CLK_noedge_posedge :	VitalDelayType := 0.530 ns;
      tpw_CLK_posedge         :	VitalDelayType := 0.660 ns;
      tperiod_CLK_posedge             :	VitalDelayType := 1.320 ns;
      trecovery_S_CLK_posedge_posedge :	VitalDelayType := 0.000 ns;---0.330 ns;
      thold_S_CLK_posedge_posedge    :	VitalDelayType := 0.530 ns;
      ticd_CLK                       :	VitalDelayType := 0.000 ns;
      tisd_D_CLK                     :	VitalDelayType := 0.000 ns;
      tisd_S_CLK                     :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of RIS : entity is TRUE;
end RIS;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library VF1;
architecture VITAL_VF of RIS is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL D_CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL S_CLK_dly	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (S_ipd, S, tipd_S);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   VitalSignalDelay (CLK_dly, CLK_ipd, ticd_CLK);
   VitalSignalDelay (D_CLK_dly, D_ipd, tisd_D_CLK);
   VitalSignalDelay (S_CLK_dly, S_ipd, tisd_S_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (CLK_dly, D_CLK_dly, S_CLK_dly)

   -- timing check results
   VARIABLE Tviol_D_CLK_S_EQ_1_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_S_EQ_1_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK_S_EQ_1	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK_S_EQ_1	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 3);
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_S_EQ_1_posedge,
          TimingData              => Tmkr_D_CLK_S_EQ_1_posedge,
          TestSignal              => D_CLK_dly,
          TestSignalName          => "D",
          TestDelay               => tisd_D_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          SetupHigh               => tsetup_D_CLK_noedge_posedge,
          SetupLow                => tsetup_D_CLK_noedge_posedge,
          HoldHigh                => thold_D_CLK_noedge_posedge,
          HoldLow                 => thold_D_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(S_CLK_dly) = '0',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/RIS",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_S_CLK_posedge,
          TimingData              => Tmkr_S_CLK_posedge,
          TestSignal              => S_CLK_dly,
          TestSignalName          => "S",
          TestDelay               => tisd_S_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          Recovery                => trecovery_S_CLK_posedge_posedge,
          Removal                 => thold_S_CLK_posedge_posedge,
          ActiveLow               => FALSE,
          CheckEnabled            => TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/RIS",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK_S_EQ_1,
          PeriodData              => PInfo_CLK_S_EQ_1,
          TestSignal              => CLK_dly,
          TestSignalName          => "CLK",
          TestDelay               => ticd_CLK,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TO_X01((S_CLK_dly) ) = '0',
          HeaderMsg               => InstancePath & "/RIS",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_S_EQ_1_posedge or Tviol_S_CLK_posedge or Pviol_CLK_S_EQ_1;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => dfftab,
        DataIn => (
               D_CLK_dly, CLK_dly, '1',NOT(S_CLK_dly)));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (S_CLK_dly'last_event, tpd_S_Q, TRUE),
                 1 => (CLK_dly'last_event, tpd_CLK_Q, TRUE)),
       Mode => VitalInertial,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;

configuration CFG_RIS_VITAL of RIS is 
        for VITAL_VF
        end for; 
end CFG_RIS_VITAL;
---------------------------------------------------------------------------------
-- VITAL model for cell ROLI
---------------------------------------------------------------------------------
LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.VITAL_timing.all;
USE IEEE.VITAL_primitives.all;
LIBRARY VF1;
USE VF1.VLOGTOVITAL_TABLES.all;

-----------------------------------------------------------------------------
--ENTITY DECLARATION
-----------------------------------------------------------------------------
ENTITY ROLI IS

GENERIC (
	tipd_IO			 : VITALDELAYTYPE01Z 	 := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
	tipd_D			 : VITALDELAYTYPE01Z 	 := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
	tipd_CLK		 : VITALDELAYTYPE01Z 	 := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
	tipd_LAT		 : VITALDELAYTYPE01Z 	 := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
	tipd_OE			 : VITALDELAYTYPE01Z 	 := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
	TimingChecksOn           : BOOLEAN               := TRUE;
	ticd_CLK		 : VITALDELAYTYPE 	 := 0 ns;
	tisd_D_CLK		 : VITALDELAYTYPE 	 := 0 ns;
	Xon                      : BOOLEAN               := TRUE;
	InstancePath             : STRING                := "*";
	MsgOn                    : BOOLEAN               := TRUE;
	tsetup_D_CLK_noedge_posedge : VITALDELAYTYPE 	 := 0.36 ns;
	thold_D_CLK_noedge_posedge : VITALDELAYTYPE 	 := 0.56 ns;
	tpw_CLK_posedge 	: VITALDELAYTYPE 	 := 0.72 ns;
	tpw_CLK_negedge 	: VITALDELAYTYPE 	 := 0 ns;
	tperiod_CLK_posedge 	: VITALDELAYTYPE 	 := 1.44 ns;
	ticd_LAT		 : VITALDELAYTYPE 	 := 0 ns;
	tisd_IO_LAT		 : VITALDELAYTYPE 	 := 0 ns;
	tsetup_IO_LAT_noedge_negedge : VITALDELAYTYPE 	 := -0.33 ns;
	thold_IO_LAT_noedge_negedge : VITALDELAYTYPE 	 := 0.53 ns;
	tpw_LAT_posedge		 : VITALDELAYTYPE 	 := 0.66 ns;
	tpw_LAT_negedge		 : VITALDELAYTYPE 	 := 0 ns;
	tperiod_LAT_posedge	 : VITALDELAYTYPE 	 := 1.32 ns;
	tpd_OE_IO		 : VITALDELAYTYPE01Z 	 := (0.64 ns, 0.64 ns, 0.64 ns, 0.64 ns, 0.64 ns, 0.64 ns);
	tpd_IO_O		 : VITALDELAYTYPE01 	 := (0.4 ns, 0.4 ns);
	tpd_CLK_O		 : VITALDELAYTYPE01 	 := (3.14 ns, 3.14 ns);
	tpd_CLK_IO		 : VITALDELAYTYPE01Z 	 := (2.74 ns, 2.74 ns,2.74 ns,2.74 ns,2.74 ns,2.74 ns);
	tpd_LAT_Q		 : VITALDELAYTYPE01 	 := (1.23 ns, 1.23 ns);
	tpd_IO_Q		 : VITALDELAYTYPE01 	 := (1.23 ns, 1.23 ns)
	);

PORT    (
	O			 : OUT   std_logic;
	Q			 : OUT   std_logic;
	IO			 : INOUT std_logic := 'U';
	D			 : IN    std_logic := 'U';
	CLK			 : IN    std_logic := 'U';
	LAT			 : IN    std_logic := 'U';
	OE			 : IN    std_logic := 'U'
	);

ATTRIBUTE VITAL_LEVEL0 OF ROLI : ENTITY IS TRUE ;

END ROLI;
-----------------------------------------------------------------------------
-- ARCHITECTURE declaration
-----------------------------------------------------------------------------
ARCHITECTURE VITAL_VF OF ROLI  IS
	ATTRIBUTE VITAL_LEVEL1 OF VITAL_VF : ARCHITECTURE IS TRUE;

	SIGNAL	IO_ipd			 : std_ulogic        := 'X';
	SIGNAL	D_ipd			 : std_ulogic        := 'X';
	SIGNAL	CLK_ipd			 : std_ulogic        := 'X';
	SIGNAL	LAT_ipd			 : std_ulogic        := 'X';
	SIGNAL	OE_ipd			 : std_ulogic        := 'X';
	SIGNAL	CLK_dly			 : std_ulogic        := 'X';
	SIGNAL	D_dly			 : std_ulogic        := 'X';
	SIGNAL	LAT_dly			 : std_ulogic        := 'X';
	SIGNAL	IO_dly			 : std_ulogic        := 'X';
BEGIN
-----------------------------------------------------------------------------
-- INPUT PATH DELAYs
-----------------------------------------------------------------------------
WIREDELAY : BLOCK
BEGIN
	VitalWireDelay( IO_ipd, IO, tipd_IO );
	VitalWireDelay( D_ipd, D, tipd_D );
	VitalWireDelay( CLK_ipd, CLK, tipd_CLK );
	VitalWireDelay( LAT_ipd, LAT, tipd_LAT );
	VitalWireDelay( OE_ipd, OE, tipd_OE );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
	VitalSignalDelay ( CLK_dly, CLK_ipd, ticd_CLK);
	VitalSignalDelay ( D_dly, D_ipd, tisd_D_CLK);
	VitalSignalDelay ( LAT_dly, LAT_ipd, ticd_LAT);
	VitalSignalDelay ( IO_dly, IO_ipd, tisd_IO_LAT);
END BLOCK;

-----------------------------------------------------------------------------
-- Behavior Section
-----------------------------------------------------------------------------
VitalBehaviour_1 : PROCESS(OE_ipd,D_dly,CLK_dly,IO_dly,LAT_dly)

VARIABLE 	Tviol_CLK_D_flag1	 : std_ulogic		 := '0';
VARIABLE 	TimingData_D_CLK1	 : VitalTimingDataType	 := VitalTimingDataInit;
VARIABLE 	Tviol_CLK_flag2		 : std_ulogic		 := '0';
VARIABLE 	PeriodData_CLK2		 : VitalPeriodDataType	 := VitalPeriodDataInit;
VARIABLE 	Tviol_CLK_flag3		 : std_ulogic		 := '0';
VARIABLE 	PeriodData_CLK3		 : VitalPeriodDataType	 := VitalPeriodDataInit;
VARIABLE 	Tviol_LAT_IO_flag4	 : std_ulogic		 := '0';
VARIABLE 	TimingData_IO_LAT4	 : VitalTimingDataType	 := VitalTimingDataInit;
VARIABLE 	Tviol_LAT_flag5		 : std_ulogic		 := '0';
VARIABLE 	PeriodData_LAT5		 : VitalPeriodDataType	 := VitalPeriodDataInit;
VARIABLE 	Tviol_LAT_flag6		 : std_ulogic		 := '0';
VARIABLE 	PeriodData_LAT6		 : VitalPeriodDataType	 := VitalPeriodDataInit;
VARIABLE 	Q_int_zd		 : std_ulogic;
VARIABLE 	VCC_zd			 : std_ulogic;
VARIABLE 	PrevDataIn0		 : std_logic_vector (0 to 3) ;
VARIABLE 	Q_zd			 : std_ulogic;
VARIABLE 	PrevDataIn1		 : std_logic_vector (0 to 3) ;
VARIABLE 	IO_zd			 : std_ulogic;
VARIABLE 	O_zd			 : std_ulogic;
VARIABLE 	OGLITCH_DATA		 : VitalGlitchDataType;
VARIABLE 	QGLITCH_DATA		 : VitalGlitchDataType;
VARIABLE 	IOGLITCH_DATA		 : VitalGlitchDataType;
VARIABLE 	Violation_Flag		 : std_ulogic;


BEGIN

--Timing Check Section

IF(TimingChecksOn) THEN
VitalSetupHoldCheck(Violation => Tviol_CLK_D_flag1,
TimingData => TimingData_D_CLK1,
TestSignal => D_dly,
TestSignalName => "D",
TestDelay => tisd_D_CLK,
RefSignal => CLK_dly,
RefSignalName => "CLK",
RefDelay => ticd_CLK,
SetupHigh => tsetup_D_CLK_noedge_posedge,
SetupLow => tsetup_D_CLK_noedge_posedge,
HoldHigh => thold_D_CLK_noedge_posedge,
HoldLow => thold_D_CLK_noedge_posedge,
CheckEnabled => ( To_X01( OE_ipd )= '1' ),
RefTransition => '/',
HeaderMsg => InstancePath & "/ROLI",
Xon => Xon,
MsgOn => MsgOn,
MsgSeverity => WARNING);

VitalPeriodPulseCheck(Violation => Tviol_CLK_flag2,
PeriodData => PeriodData_CLK2,
TestSignal => CLK_dly,
TestSignalName => "CLK",
TestDelay => ticd_CLK,
Period => 0 ns,
PulseWidthHigh => tpw_CLK_posedge,
PulseWidthLow => tpw_CLK_negedge,
CheckEnabled => ( To_X01( OE_ipd )= '1' ),
HeaderMsg => InstancePath & "/ROLI",
Xon => Xon,
MsgOn => MsgOn,
MsgSeverity => WARNING);

VitalPeriodPulseCheck(Violation => Tviol_CLK_flag3,
PeriodData => PeriodData_CLK3,
TestSignal => CLK_dly,
TestSignalName => "CLK",
TestDelay => ticd_CLK,
Period => tperiod_CLK_posedge,
PulseWidthHigh => 0 ns,
PulseWidthLow => 0 ns,
CheckEnabled => posedge( CLK_dly'LAST_VALUE, CLK_dly ) AND ( To_X01( OE_ipd )= '1' ),
HeaderMsg => InstancePath & "/ROLI",
Xon => Xon,
MsgOn => MsgOn,
MsgSeverity => WARNING);

VitalSetupHoldCheck(Violation => Tviol_LAT_IO_flag4,
TimingData => TimingData_IO_LAT4,
TestSignal => IO_dly,
TestSignalName => "IO",
TestDelay => tisd_IO_LAT,
RefSignal => LAT_dly,
RefSignalName => "LAT",
RefDelay => ticd_LAT,
SetupHigh => tsetup_IO_LAT_noedge_negedge,
SetupLow => tsetup_IO_LAT_noedge_negedge,
HoldHigh => thold_IO_LAT_noedge_negedge,
HoldLow => thold_IO_LAT_noedge_negedge,
CheckEnabled => TRUE,
RefTransition => '\',
HeaderMsg => InstancePath & "/ROLI",
Xon => Xon,
MsgOn => MsgOn,
MsgSeverity => WARNING);

VitalPeriodPulseCheck(Violation => Tviol_LAT_flag5,
PeriodData => PeriodData_LAT5,
TestSignal => LAT_dly,
TestSignalName => "LAT",
TestDelay => ticd_LAT,
Period => 0 ns,
PulseWidthHigh => tpw_LAT_posedge,
PulseWidthLow => tpw_LAT_negedge,
CheckEnabled => TRUE,
HeaderMsg => InstancePath & "/ROLI",
Xon => Xon,
MsgOn => MsgOn,
MsgSeverity => WARNING);

VitalPeriodPulseCheck(Violation => Tviol_LAT_flag6,
PeriodData => PeriodData_LAT6,
TestSignal => LAT_dly,
TestSignalName => "LAT",
TestDelay => ticd_LAT,
Period => tperiod_LAT_posedge,
PulseWidthHigh => 0 ns,
PulseWidthLow => 0 ns,
CheckEnabled => posedge( LAT_dly'LAST_VALUE, LAT_dly ),
HeaderMsg => InstancePath & "/ROLI",
Xon => Xon,
MsgOn => MsgOn,
MsgSeverity => WARNING);

END IF;   -- Timing Check Section

--Functionality Section

Violation_Flag	 := (((((Tviol_CLK_D_flag1 or Tviol_CLK_flag2) or Tviol_CLK_flag3) or Tviol_LAT_IO_flag4) or Tviol_LAT_flag5) or Tviol_LAT_flag6);
VCC_zd		 := '1';
VitalStateTable(
StateTable => dfftab,
DataIn => std_logic_vector'(D_dly,CLK_dly,VCC_zd,VCC_zd),
Result => Q_int_zd	,
PreviousDataIn => PrevDataIn0);
Q_int_zd	 := (Violation_Flag xor Q_int_zd);

IO_zd		 := VitalBUFIF1(Q_int_zd,OE_ipd);
O_zd		 := VitalBUF(IO_dly);

VitalStateTable(
StateTable => latchtab,
DataIn => std_logic_vector'(IO_dly,LAT_dly,VCC_zd,VCC_zd),
Result => Q_zd		,
PreviousDataIn => PrevDataIn1);
Q_zd		 := (Violation_Flag xor Q_zd);


--PathDelay Section

 VitalPathDelay01 ( O, OGLITCH_DATA, "O", O_zd,
	Paths => (
	0 => ( IO_dly'LAST_EVENT, tpd_IO_O, TRUE ),
	1 => ( CLK_dly'LAST_EVENT, tpd_CLK_O, TRUE ) ),
	DefaultDelay=>VitalZeroDelay01,
	Mode=>VitalInertial,
	XON=>TRUE,
	MsgOn=>TRUE,
	MsgSeverity=>WARNING );

 VitalPathDelay01 ( Q, QGLITCH_DATA, "Q", Q_zd,
	Paths => (
	0 => ( LAT_dly'LAST_EVENT, tpd_LAT_Q, TRUE ),
	1 => ( IO_dly'LAST_EVENT, tpd_IO_Q, TRUE ) ),
	DefaultDelay=>VitalZeroDelay01,
	Mode=>VitalInertial,
	XON=>TRUE,
	MsgOn=>TRUE,
	MsgSeverity=>WARNING );

 VitalPathDelay01Z ( IO, IOGLITCH_DATA, "IO", IO_zd,
	Paths => (
	0 => ( OE_ipd'LAST_EVENT, tpd_OE_IO, TRUE ),
	1 => ( CLK_dly'LAST_EVENT, tpd_CLK_IO, TRUE ) ),
	DefaultDelay=>VitalZeroDelay01Z,
	Mode=>VitalInertial,
	XON=>TRUE,
	MsgOn=>TRUE,
	MsgSeverity=>WARNING );


END PROCESS VitalBehaviour_1;
END VITAL_VF;
configuration CFG_ROLI_VITAL of ROLI is 
        for VITAL_VF
        end for; 
end CFG_ROLI_VITAL;
---------------------------------------------------------------------------------
-- VITAL model for cell ROLIR
---------------------------------------------------------------------------------
LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.VITAL_timing.all;
USE IEEE.VITAL_primitives.all;
LIBRARY VF1;
USE VF1.VLOGTOVITAL_TABLES.all;

-----------------------------------------------------------------------------
--ENTITY DECLARATION
-----------------------------------------------------------------------------
ENTITY ROLIR IS

GENERIC (
	tipd_IO			 : VITALDELAYTYPE01Z 	 := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
	tipd_D			 : VITALDELAYTYPE01Z 	 := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
	tipd_CLK		 : VITALDELAYTYPE01Z 	 := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
	tipd_LAT		 : VITALDELAYTYPE01Z 	 := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
	tipd_OE			 : VITALDELAYTYPE01Z 	 := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
	tipd_R			 : VITALDELAYTYPE01Z 	 := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
	TimingChecksOn           : BOOLEAN               := TRUE;
	ticd_CLK		 : VITALDELAYTYPE 	 := 0 ns;
	tisd_D_CLK		 : VITALDELAYTYPE 	 := 0 ns;
	Xon                      : BOOLEAN               := TRUE;
	InstancePath             : STRING                := "*";
	MsgOn                    : BOOLEAN               := TRUE;
	tsetup_D_CLK_noedge_posedge : VITALDELAYTYPE 	 := 0.36 ns;
	thold_D_CLK_noedge_posedge : VITALDELAYTYPE 	 := 0.56 ns;
	tpw_CLK_posedge 	: VITALDELAYTYPE 	 := 0.72 ns;
	tpw_CLK_negedge 	: VITALDELAYTYPE 	 := 0 ns;
	tperiod_CLK_posedge 	: VITALDELAYTYPE 	 := 1.44 ns;
        trecovery_R_CLK_posedge_posedge : VitalDelayType := 0.330 ns;
        thold_R_CLK_posedge_posedge :     VitalDelayType := 0.530 ns;
	ticd_LAT		 : VITALDELAYTYPE 	 := 0 ns;
	tisd_IO_LAT		 : VITALDELAYTYPE 	 := 0 ns;
        tisd_R_CLK                     :  VitalDelayType := 0.000 ns;
	tsetup_IO_LAT_noedge_negedge : VITALDELAYTYPE 	 := 0.33 ns;
	thold_IO_LAT_noedge_negedge : VITALDELAYTYPE 	 := 0.53 ns;
	tpw_LAT_posedge		 : VITALDELAYTYPE 	 := 0.66 ns;
	tpw_LAT_negedge		 : VITALDELAYTYPE 	 := 0 ns;
	tperiod_LAT_posedge	 : VITALDELAYTYPE 	 := 1.32 ns;
	tpd_OE_IO		 : VITALDELAYTYPE01Z 	 := (0.64 ns, 0.64 ns, 0.64 ns, 0.64 ns, 0.64 ns, 0.64 ns);
	tpd_IO_O		 : VITALDELAYTYPE01 	 := (0.4 ns, 0.4 ns);
	tpd_CLK_O		 : VITALDELAYTYPE01 	 := (3.14 ns, 3.14 ns);
        tpd_CLK_IO               : VITALDELAYTYPE01Z     := (2.74 ns, 2.74 ns,2.74 ns,2.74 ns,2.74 ns,2.74 ns);
	tpd_R_O		         : VITALDELAYTYPE01 	 := (3.14 ns, 3.14 ns);
        tpd_R_IO                 : VitalDelayType01Z      := (2.74 ns, 2.74 ns,2.74 ns, 2.74 ns,2.74 ns,2.74 ns);
	tpd_LAT_Q		 : VITALDELAYTYPE01 	 := (1.23 ns, 1.23 ns);
	tpd_IO_Q		 : VITALDELAYTYPE01 	 := (1.23 ns, 1.23 ns)
	);

PORT    (
	O			 : OUT   std_logic;
	Q			 : OUT   std_logic;
	IO			 : INOUT std_logic := 'U';
	D			 : IN    std_logic := 'U';
	CLK			 : IN    std_logic := 'U';
	LAT			 : IN    std_logic := 'U';
	OE			 : IN    std_logic := 'U';
        R                        : IN    std_logic:= 'U'
	);

ATTRIBUTE VITAL_LEVEL0 OF ROLIR : ENTITY IS TRUE ;

END ROLIR;
-----------------------------------------------------------------------------
-- ARCHITECTURE declaration
-----------------------------------------------------------------------------
ARCHITECTURE VITAL_VF OF ROLIR  IS
	ATTRIBUTE VITAL_LEVEL1 OF VITAL_VF : ARCHITECTURE IS TRUE;

	SIGNAL	IO_ipd			 : std_ulogic        := 'X';
	SIGNAL	D_ipd			 : std_ulogic        := 'X';
	SIGNAL	CLK_ipd			 : std_ulogic        := 'X';
	SIGNAL	LAT_ipd			 : std_ulogic        := 'X';
	SIGNAL	OE_ipd			 : std_ulogic        := 'X';
        SIGNAL  R_ipd                    : std_ulogic        := 'X';
	SIGNAL	CLK_dly			 : std_ulogic        := 'X';
	SIGNAL	D_dly			 : std_ulogic        := 'X';
	SIGNAL	LAT_dly			 : std_ulogic        := 'X';
	SIGNAL	IO_dly			 : std_ulogic        := 'X';
        SIGNAL  R_CLK_dly                : std_ulogic        := 'X';

BEGIN
-----------------------------------------------------------------------------
-- INPUT PATH DELAYs
-----------------------------------------------------------------------------
WIREDELAY : BLOCK
BEGIN
	VitalWireDelay( IO_ipd, IO, tipd_IO );
	VitalWireDelay( D_ipd, D, tipd_D );
	VitalWireDelay( CLK_ipd, CLK, tipd_CLK );
	VitalWireDelay( LAT_ipd, LAT, tipd_LAT );
	VitalWireDelay( OE_ipd, OE, tipd_OE );
        VitalWireDelay (R_ipd, R, tipd_R);

END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
	VitalSignalDelay ( CLK_dly, CLK_ipd, ticd_CLK);
	VitalSignalDelay ( D_dly, D_ipd, tisd_D_CLK);
	VitalSignalDelay ( LAT_dly, LAT_ipd, ticd_LAT);
	VitalSignalDelay ( IO_dly, IO_ipd, tisd_IO_LAT);
        VitalSignalDelay ( R_CLK_dly, R_ipd, tisd_R_CLK);

END BLOCK;

-----------------------------------------------------------------------------
-- Behavior Section
-----------------------------------------------------------------------------
VitalBehaviour_1 : PROCESS(OE_ipd,D_dly,CLK_dly,IO_dly,LAT_dly,R_CLK_dly)

VARIABLE 	Tviol_CLK_D_flag1	 : std_ulogic		 := '0';
VARIABLE 	TimingData_D_CLK1	 : VitalTimingDataType	 := VitalTimingDataInit;
VARIABLE        Tviol_R_CLK_OE_EQ_1_posedge : std_ulogic := '0';
VARIABLE        Tmkr_R_CLK_OE_EQ_1_posedge : VitalTimingDataType := VitalTimingDataInit;
VARIABLE 	Tviol_CLK_flag2		 : std_ulogic		 := '0';
VARIABLE 	PeriodData_CLK2		 : VitalPeriodDataType	 := VitalPeriodDataInit;
VARIABLE 	Tviol_CLK_flag3		 : std_ulogic		 := '0';
VARIABLE 	PeriodData_CLK3		 : VitalPeriodDataType	 := VitalPeriodDataInit;
VARIABLE 	Tviol_LAT_IO_flag4	 : std_ulogic		 := '0';
VARIABLE 	TimingData_IO_LAT4	 : VitalTimingDataType	 := VitalTimingDataInit;
VARIABLE 	Tviol_LAT_flag5		 : std_ulogic		 := '0';
VARIABLE 	PeriodData_LAT5		 : VitalPeriodDataType	 := VitalPeriodDataInit;
VARIABLE 	Tviol_LAT_flag6		 : std_ulogic		 := '0';
VARIABLE 	PeriodData_LAT6		 : VitalPeriodDataType	 := VitalPeriodDataInit;
VARIABLE 	Q_int_zd		 : std_ulogic;
VARIABLE 	VCC_zd			 : std_ulogic;
VARIABLE 	PrevDataIn0		 : std_logic_vector (0 to 3) ;
VARIABLE 	Q_zd			 : std_ulogic;
VARIABLE 	PrevDataIn1		 : std_logic_vector (0 to 3) ;
VARIABLE 	IO_zd			 : std_ulogic;
VARIABLE 	O_zd			 : std_ulogic;
VARIABLE 	OGLITCH_DATA		 : VitalGlitchDataType;
VARIABLE 	QGLITCH_DATA		 : VitalGlitchDataType;
VARIABLE 	IOGLITCH_DATA		 : VitalGlitchDataType;
VARIABLE 	Violation_Flag		 : std_ulogic;


BEGIN

--Timing Check Section

IF(TimingChecksOn) THEN
VitalSetupHoldCheck(Violation => Tviol_CLK_D_flag1,
TimingData => TimingData_D_CLK1,
TestSignal => D_dly,
TestSignalName => "D",
TestDelay => tisd_D_CLK,
RefSignal => CLK_dly,
RefSignalName => "CLK",
RefDelay => ticd_CLK,
SetupHigh => tsetup_D_CLK_noedge_posedge,
SetupLow => tsetup_D_CLK_noedge_posedge,
HoldHigh => thold_D_CLK_noedge_posedge,
HoldLow => thold_D_CLK_noedge_posedge,
CheckEnabled => ( To_X01( OE_ipd AND NOT(R_CLK_dly))= '1' ),
RefTransition => '/',
HeaderMsg => InstancePath & "/ROLIR",
Xon => Xon,
MsgOn => MsgOn,
MsgSeverity => WARNING);

VitalPeriodPulseCheck(Violation => Tviol_CLK_flag2,
PeriodData => PeriodData_CLK2,
TestSignal => CLK_dly,
TestSignalName => "CLK",
TestDelay => ticd_CLK,
Period => 0 ns,
PulseWidthHigh => tpw_CLK_posedge,
PulseWidthLow => tpw_CLK_negedge,
CheckEnabled => ( To_X01( OE_ipd AND NOT(R_CLK_dly))= '1' ),
HeaderMsg => InstancePath & "/ROLIR",
Xon => Xon,
MsgOn => MsgOn,
MsgSeverity => WARNING);

VitalPeriodPulseCheck(Violation => Tviol_CLK_flag3,
PeriodData => PeriodData_CLK3,
TestSignal => CLK_dly,
TestSignalName => "CLK",
TestDelay => ticd_CLK,
Period => tperiod_CLK_posedge,
PulseWidthHigh => 0 ns,
PulseWidthLow => 0 ns,
CheckEnabled => posedge( CLK_dly'LAST_VALUE, CLK_dly ) AND ( To_X01( OE_ipd AND NOT(R_CLK_dly))= '1' ),
HeaderMsg => InstancePath & "/ROLIR",
Xon => Xon,
MsgOn => MsgOn,
MsgSeverity => WARNING);

VitalSetupHoldCheck(Violation => Tviol_LAT_IO_flag4,
TimingData => TimingData_IO_LAT4,
TestSignal => IO_dly,
TestSignalName => "IO",
TestDelay => tisd_IO_LAT,
RefSignal => LAT_dly,
RefSignalName => "LAT",
RefDelay => ticd_LAT,
SetupHigh => tsetup_IO_LAT_noedge_negedge,
SetupLow => tsetup_IO_LAT_noedge_negedge,
HoldHigh => thold_IO_LAT_noedge_negedge,
HoldLow => thold_IO_LAT_noedge_negedge,
CheckEnabled => TRUE,
RefTransition => '\',
HeaderMsg => InstancePath & "/ROLIR",
Xon => Xon,
MsgOn => MsgOn,
MsgSeverity => WARNING);

VitalPeriodPulseCheck(Violation => Tviol_LAT_flag5,
PeriodData => PeriodData_LAT5,
TestSignal => LAT_dly,
TestSignalName => "LAT",
TestDelay => ticd_LAT,
Period => 0 ns,
PulseWidthHigh => tpw_LAT_posedge,
PulseWidthLow => tpw_LAT_negedge,
CheckEnabled => TRUE,
HeaderMsg => InstancePath & "/ROLIR",
Xon => Xon,
MsgOn => MsgOn,
MsgSeverity => WARNING);

VitalPeriodPulseCheck(Violation => Tviol_LAT_flag6,
PeriodData => PeriodData_LAT6,
TestSignal => LAT_dly,
TestSignalName => "LAT",
TestDelay => ticd_LAT,
Period => tperiod_LAT_posedge,
PulseWidthHigh => 0 ns,
PulseWidthLow => 0 ns,
CheckEnabled => posedge( LAT_dly'LAST_VALUE, LAT_dly ),
HeaderMsg => InstancePath & "/ROLIR",
Xon => Xon,
MsgOn => MsgOn,
MsgSeverity => WARNING);

VitalRecoveryRemovalCheck ( Violation  => Tviol_R_CLK_OE_EQ_1_posedge,
TimingData  => Tmkr_R_CLK_OE_EQ_1_posedge,
TestSignal  => R_CLK_dly,
TestSignalName  => "R",
TestDelay  => tisd_R_CLK,
RefSignal  => CLK_dly,
RefSignalName  => "CLK",
RefDelay  => ticd_CLK,
Recovery  => trecovery_R_CLK_posedge_posedge,
Removal   => thold_R_CLK_posedge_posedge,
ActiveLow  => FALSE,
CheckEnabled  => TO_X01(OE_ipd) = '1',
RefTransition  => 'R',
HeaderMsg  => InstancePath & "/ROLIR",
Xon  => Xon,
MsgOn  => MsgOn,
MsgSeverity  => WARNING);


END IF;   -- Timing Check Section

--Functionality Section

Violation_Flag	 := Tviol_CLK_D_flag1 or Tviol_CLK_flag2 or Tviol_CLK_flag3 or Tviol_LAT_IO_flag4 or Tviol_LAT_flag5 or Tviol_LAT_flag6 or Tviol_R_CLK_OE_EQ_1_posedge;
VCC_zd		 := '1';
VitalStateTable(
StateTable => dfftab,
DataIn => std_logic_vector'(D_dly,CLK_dly,NOT(R_CLK_dly),VCC_zd),
Result => Q_int_zd	,
PreviousDataIn => PrevDataIn0);
Q_int_zd	 := (Violation_Flag xor Q_int_zd);

IO_zd		 := VitalBUFIF1(Q_int_zd,OE_ipd);
O_zd		 := VitalBUF(IO_dly);

VitalStateTable(
StateTable => latchtab,
DataIn => std_logic_vector'(IO_dly,LAT_dly,VCC_zd,VCC_zd),
Result => Q_zd		,
PreviousDataIn => PrevDataIn1);
--Q_zd		 := (Violation_Flag xor Q_zd);


--PathDelay Section

 VitalPathDelay01 ( O, OGLITCH_DATA, "O", O_zd,
	Paths => (
	0 => ( IO_dly'LAST_EVENT, tpd_IO_O, TRUE ),
	1 => ( CLK_dly'LAST_EVENT, tpd_CLK_O, TRUE ),
        2 => ( R_CLK_dly'LAST_EVENT, tpd_R_O, TRUE)),
	DefaultDelay=>VitalZeroDelay01,
	Mode=>VitalInertial,
	XON=>TRUE,
	MsgOn=>TRUE,
	MsgSeverity=>WARNING );

 VitalPathDelay01 ( Q, QGLITCH_DATA, "Q", Q_zd,
	Paths => (
	0 => ( LAT_dly'LAST_EVENT, tpd_LAT_Q, TRUE ),
	1 => ( IO_dly'LAST_EVENT, tpd_IO_Q, TRUE ) ),
	DefaultDelay=>VitalZeroDelay01,
	Mode=>VitalInertial,
	XON=>TRUE,
	MsgOn=>TRUE,
	MsgSeverity=>WARNING );

 VitalPathDelay01Z ( IO, IOGLITCH_DATA, "IO", IO_zd,
	Paths => (
	0 => ( OE_ipd'LAST_EVENT, tpd_OE_IO, TRUE ),
        1 => ( CLK_dly'LAST_EVENT, tpd_CLK_IO, TRUE ),
        2 => ( R_CLK_dly'LAST_EVENT, tpd_R_IO, TRUE ) ),
	DefaultDelay=>VitalZeroDelay01Z,
	Mode=>VitalInertial,
	XON=>TRUE,
	MsgOn=>TRUE,
	MsgSeverity=>WARNING );


END PROCESS VitalBehaviour_1;
END VITAL_VF;
configuration CFG_ROLIR_VITAL of ROLIR is 
        for VITAL_VF
        end for; 
end CFG_ROLIR_VITAL;
---------------------------------------------------------------------------------
-- VITAL model for cell ROLIS
---------------------------------------------------------------------------------
LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.VITAL_timing.all;
USE IEEE.VITAL_primitives.all;
LIBRARY VF1;
USE VF1.VLOGTOVITAL_TABLES.all;

-----------------------------------------------------------------------------
--ENTITY DECLARATION
-----------------------------------------------------------------------------
ENTITY ROLIS IS

GENERIC (
	tipd_IO			 : VITALDELAYTYPE01Z 	 := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
	tipd_D			 : VITALDELAYTYPE01Z 	 := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
	tipd_CLK		 : VITALDELAYTYPE01Z 	 := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
	tipd_LAT		 : VITALDELAYTYPE01Z 	 := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
	tipd_OE			 : VITALDELAYTYPE01Z 	 := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
	tipd_S			 : VITALDELAYTYPE01Z 	 := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
	TimingChecksOn           : BOOLEAN               := TRUE;
	ticd_CLK		 : VITALDELAYTYPE 	 := 0 ns;
	tisd_D_CLK		 : VITALDELAYTYPE 	 := 0 ns;
	Xon                      : BOOLEAN               := TRUE;
	InstancePath             : STRING                := "*";
	MsgOn                    : BOOLEAN               := TRUE;
	tsetup_D_CLK_noedge_posedge : VITALDELAYTYPE 	 := 0.36 ns;
	thold_D_CLK_noedge_posedge : VITALDELAYTYPE 	 := 0.56 ns;
	tpw_CLK_posedge 	: VITALDELAYTYPE 	 := 0.72 ns;
	tpw_CLK_negedge 	: VITALDELAYTYPE 	 := 0 ns;
	tperiod_CLK_posedge 	: VITALDELAYTYPE 	 := 1.44 ns;
        trecovery_S_CLK_posedge_posedge : VitalDelayType := 0.330 ns;
        thold_S_CLK_posedge_posedge :     VitalDelayType := 0.530 ns;
	ticd_LAT		 : VITALDELAYTYPE 	 := 0 ns;
	tisd_IO_LAT		 : VITALDELAYTYPE 	 := 0 ns;
        tisd_S_CLK                     :  VitalDelayType := 0.000 ns;
	tsetup_IO_LAT_noedge_negedge : VITALDELAYTYPE 	 := 0.33 ns;
	thold_IO_LAT_noedge_negedge : VITALDELAYTYPE 	 := 0.53 ns;
	tpw_LAT_posedge		 : VITALDELAYTYPE 	 := 0.66 ns;
	tpw_LAT_negedge		 : VITALDELAYTYPE 	 := 0 ns;
	tperiod_LAT_posedge	 : VITALDELAYTYPE 	 := 1.32 ns;
	tpd_OE_IO		 : VITALDELAYTYPE01Z 	 := (0.64 ns, 0.64 ns, 0.64 ns, 0.64 ns, 0.64 ns, 0.64 ns);
	tpd_IO_O		 : VITALDELAYTYPE01 	 := (0.4 ns, 0.4 ns);
	tpd_CLK_O		 : VITALDELAYTYPE01 	 := (3.14 ns, 3.14 ns);
        tpd_CLK_IO               : VITALDELAYTYPE01Z     := (2.74 ns, 2.74 ns,2.74 ns,2.74 ns,2.74 ns,2.74 ns);
	tpd_S_O		         : VITALDELAYTYPE01 	 := (3.14 ns, 3.14 ns);
        tpd_S_IO                 : VitalDelayType01Z      := (2.74 ns, 2.74 ns,2.74 ns, 2.74 ns,2.74 ns,2.74 ns);
	tpd_LAT_Q		 : VITALDELAYTYPE01 	 := (1.23 ns, 1.23 ns);
	tpd_IO_Q		 : VITALDELAYTYPE01 	 := (1.23 ns, 1.23 ns)
	);

PORT    (
	O			 : OUT   std_logic;
	Q			 : OUT   std_logic;
	IO			 : INOUT std_logic := 'U';
	D			 : IN    std_logic := 'U';
	CLK			 : IN    std_logic := 'U';
	LAT			 : IN    std_logic := 'U';
	OE			 : IN    std_logic := 'U';
        S                        : IN    std_logic:= 'U'
	);

ATTRIBUTE VITAL_LEVEL0 OF ROLIS : ENTITY IS TRUE ;

END ROLIS;
-----------------------------------------------------------------------------
-- ARCHITECTURE declaration
-----------------------------------------------------------------------------
ARCHITECTURE VITAL_VF OF ROLIS  IS
	ATTRIBUTE VITAL_LEVEL1 OF VITAL_VF : ARCHITECTURE IS TRUE;

	SIGNAL	IO_ipd			 : std_ulogic        := 'X';
	SIGNAL	D_ipd			 : std_ulogic        := 'X';
	SIGNAL	CLK_ipd			 : std_ulogic        := 'X';
	SIGNAL	LAT_ipd			 : std_ulogic        := 'X';
	SIGNAL	OE_ipd			 : std_ulogic        := 'X';
        SIGNAL  S_ipd                    : std_ulogic        := 'X';
	SIGNAL	CLK_dly			 : std_ulogic        := 'X';
	SIGNAL	D_dly			 : std_ulogic        := 'X';
	SIGNAL	LAT_dly			 : std_ulogic        := 'X';
	SIGNAL	IO_dly			 : std_ulogic        := 'X';
        SIGNAL  S_CLK_dly                : std_ulogic        := 'X';

BEGIN
-----------------------------------------------------------------------------
-- INPUT PATH DELAYs
-----------------------------------------------------------------------------
WIREDELAY : BLOCK
BEGIN
	VitalWireDelay( IO_ipd, IO, tipd_IO );
	VitalWireDelay( D_ipd, D, tipd_D );
	VitalWireDelay( CLK_ipd, CLK, tipd_CLK );
	VitalWireDelay( LAT_ipd, LAT, tipd_LAT );
	VitalWireDelay( OE_ipd, OE, tipd_OE );
        VitalWireDelay( S_ipd, S, tipd_S);

END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
	VitalSignalDelay ( CLK_dly, CLK_ipd, ticd_CLK);
	VitalSignalDelay ( D_dly, D_ipd, tisd_D_CLK);
	VitalSignalDelay ( LAT_dly, LAT_ipd, ticd_LAT);
	VitalSignalDelay ( IO_dly, IO_ipd, tisd_IO_LAT);
        VitalSignalDelay ( S_CLK_dly, S_ipd, tisd_S_CLK);

END BLOCK;

-----------------------------------------------------------------------------
-- Behavior Section
-----------------------------------------------------------------------------
VitalBehaviour_1 : PROCESS(OE_ipd,D_dly,CLK_dly,IO_dly,LAT_dly,S_CLK_dly)

VARIABLE 	Tviol_CLK_D_flag1	 : std_ulogic		 := '0';
VARIABLE 	TimingData_D_CLK1	 : VitalTimingDataType	 := VitalTimingDataInit;
VARIABLE        Tviol_S_CLK_OE_EQ_1_posedge : std_ulogic := '0';
VARIABLE        Tmkr_S_CLK_OE_EQ_1_posedge : VitalTimingDataType := VitalTimingDataInit;
VARIABLE 	Tviol_CLK_flag2		 : std_ulogic		 := '0';
VARIABLE 	PeriodData_CLK2		 : VitalPeriodDataType	 := VitalPeriodDataInit;
VARIABLE 	Tviol_CLK_flag3		 : std_ulogic		 := '0';
VARIABLE 	PeriodData_CLK3		 : VitalPeriodDataType	 := VitalPeriodDataInit;
VARIABLE 	Tviol_LAT_IO_flag4	 : std_ulogic		 := '0';
VARIABLE 	TimingData_IO_LAT4	 : VitalTimingDataType	 := VitalTimingDataInit;
VARIABLE 	Tviol_LAT_flag5		 : std_ulogic		 := '0';
VARIABLE 	PeriodData_LAT5		 : VitalPeriodDataType	 := VitalPeriodDataInit;
VARIABLE 	Tviol_LAT_flag6		 : std_ulogic		 := '0';
VARIABLE 	PeriodData_LAT6		 : VitalPeriodDataType	 := VitalPeriodDataInit;
VARIABLE 	Q_int_zd		 : std_ulogic;
VARIABLE 	VCC_zd			 : std_ulogic;
VARIABLE 	PrevDataIn0		 : std_logic_vector (0 to 3) ;
VARIABLE 	Q_zd			 : std_ulogic;
VARIABLE 	PrevDataIn1		 : std_logic_vector (0 to 3) ;
VARIABLE 	IO_zd			 : std_ulogic;
VARIABLE 	O_zd			 : std_ulogic;
VARIABLE 	OGLITCH_DATA		 : VitalGlitchDataType;
VARIABLE 	QGLITCH_DATA		 : VitalGlitchDataType;
VARIABLE 	IOGLITCH_DATA		 : VitalGlitchDataType;
VARIABLE 	Violation_Flag		 : std_ulogic;


BEGIN

--Timing Check Section

IF(TimingChecksOn) THEN
VitalSetupHoldCheck(Violation => Tviol_CLK_D_flag1,
TimingData => TimingData_D_CLK1,
TestSignal => D_dly,
TestSignalName => "D",
TestDelay => tisd_D_CLK,
RefSignal => CLK_dly,
RefSignalName => "CLK",
RefDelay => ticd_CLK,
SetupHigh => tsetup_D_CLK_noedge_posedge,
SetupLow => tsetup_D_CLK_noedge_posedge,
HoldHigh => thold_D_CLK_noedge_posedge,
HoldLow => thold_D_CLK_noedge_posedge,
CheckEnabled => ( To_X01( OE_ipd AND NOT(S_CLK_dly))= '1' ),
RefTransition => '/',
HeaderMsg => InstancePath & "/ROLIS",
Xon => Xon,
MsgOn => MsgOn,
MsgSeverity => WARNING);

VitalPeriodPulseCheck(Violation => Tviol_CLK_flag2,
PeriodData => PeriodData_CLK2,
TestSignal => CLK_dly,
TestSignalName => "CLK",
TestDelay => ticd_CLK,
Period => 0 ns,
PulseWidthHigh => tpw_CLK_posedge,
PulseWidthLow => tpw_CLK_negedge,
CheckEnabled => ( To_X01( OE_ipd AND NOT(S_CLK_dly))= '1' ),
HeaderMsg => InstancePath & "/ROLIS",
Xon => Xon,
MsgOn => MsgOn,
MsgSeverity => WARNING);

VitalPeriodPulseCheck(Violation => Tviol_CLK_flag3,
PeriodData => PeriodData_CLK3,
TestSignal => CLK_dly,
TestSignalName => "CLK",
TestDelay => ticd_CLK,
Period => tperiod_CLK_posedge,
PulseWidthHigh => 0 ns,
PulseWidthLow => 0 ns,
CheckEnabled => posedge( CLK_dly'LAST_VALUE, CLK_dly ) AND ( To_X01( OE_ipd AND NOT(S_CLK_dly))= '1' ),
HeaderMsg => InstancePath & "/ROLIS",
Xon => Xon,
MsgOn => MsgOn,
MsgSeverity => WARNING);

VitalSetupHoldCheck(Violation => Tviol_LAT_IO_flag4,
TimingData => TimingData_IO_LAT4,
TestSignal => IO_dly,
TestSignalName => "IO",
TestDelay => tisd_IO_LAT,
RefSignal => LAT_dly,
RefSignalName => "LAT",
RefDelay => ticd_LAT,
SetupHigh => tsetup_IO_LAT_noedge_negedge,
SetupLow => tsetup_IO_LAT_noedge_negedge,
HoldHigh => thold_IO_LAT_noedge_negedge,
HoldLow => thold_IO_LAT_noedge_negedge,
CheckEnabled => TRUE,
RefTransition => '\',
HeaderMsg => InstancePath & "/ROLIS",
Xon => Xon,
MsgOn => MsgOn,
MsgSeverity => WARNING);

VitalPeriodPulseCheck(Violation => Tviol_LAT_flag5,
PeriodData => PeriodData_LAT5,
TestSignal => LAT_dly,
TestSignalName => "LAT",
TestDelay => ticd_LAT,
Period => 0 ns,
PulseWidthHigh => tpw_LAT_posedge,
PulseWidthLow => tpw_LAT_negedge,
CheckEnabled => TRUE,
HeaderMsg => InstancePath & "/ROLIS",
Xon => Xon,
MsgOn => MsgOn,
MsgSeverity => WARNING);

VitalPeriodPulseCheck(Violation => Tviol_LAT_flag6,
PeriodData => PeriodData_LAT6,
TestSignal => LAT_dly,
TestSignalName => "LAT",
TestDelay => ticd_LAT,
Period => tperiod_LAT_posedge,
PulseWidthHigh => 0 ns,
PulseWidthLow => 0 ns,
CheckEnabled => posedge( LAT_dly'LAST_VALUE, LAT_dly ),
HeaderMsg => InstancePath & "/ROLIS",
Xon => Xon,
MsgOn => MsgOn,
MsgSeverity => WARNING);

VitalRecoveryRemovalCheck ( Violation  => Tviol_S_CLK_OE_EQ_1_posedge,
TimingData  => Tmkr_S_CLK_OE_EQ_1_posedge,
TestSignal  => S_CLK_dly,
TestSignalName  => "S",
TestDelay  => tisd_S_CLK,
RefSignal  => CLK_dly,
RefSignalName  => "CLK",
RefDelay  => ticd_CLK,
Recovery  => trecovery_S_CLK_posedge_posedge,
Removal   => thold_S_CLK_posedge_posedge,
ActiveLow  => FALSE,
CheckEnabled  => TO_X01(OE_ipd) = '1',
RefTransition  => 'R',
HeaderMsg  => InstancePath & "/ROLIS",
Xon  => Xon,
MsgOn  => MsgOn,
MsgSeverity  => WARNING);


END IF;   -- Timing Check Section

--Functionality Section

Violation_Flag	 := (((((Tviol_CLK_D_flag1 or Tviol_CLK_flag2) or Tviol_CLK_flag3) or Tviol_LAT_IO_flag4) or Tviol_LAT_flag5) or Tviol_LAT_flag6 or Tviol_S_CLK_OE_EQ_1_posedge);
VCC_zd		 := '1';
VitalStateTable(
StateTable => dfftab,
DataIn => std_logic_vector'(D_dly,CLK_dly,VCC_zd,NOT(S_CLK_dly)),
Result => Q_int_zd	,
PreviousDataIn => PrevDataIn0);
Q_int_zd	 := (Violation_Flag xor Q_int_zd);

IO_zd		 := VitalBUFIF1(Q_int_zd,OE_ipd);
O_zd		 := VitalBUF(IO_dly);

VitalStateTable(
StateTable => latchtab,
DataIn => std_logic_vector'(IO_dly,LAT_dly,VCC_zd,VCC_zd),
Result => Q_zd		,
PreviousDataIn => PrevDataIn1);
Q_zd		 := (Violation_Flag xor Q_zd);


--PathDelay Section

 VitalPathDelay01 ( O, OGLITCH_DATA, "O", O_zd,
	Paths => (
	0 => ( IO_dly'LAST_EVENT, tpd_IO_O, TRUE ),
	1 => ( CLK_dly'LAST_EVENT, tpd_CLK_O, TRUE ),
        2 =>  (S_CLK_dly'LAST_EVENT, tpd_S_O, TRUE)),
	DefaultDelay=>VitalZeroDelay01,
	Mode=>VitalInertial,
	XON=>TRUE,
	MsgOn=>TRUE,
	MsgSeverity=>WARNING );

 VitalPathDelay01 ( Q, QGLITCH_DATA, "Q", Q_zd,
	Paths => (
	0 => ( LAT_dly'LAST_EVENT, tpd_LAT_Q, TRUE ),
	1 => ( IO_dly'LAST_EVENT, tpd_IO_Q, TRUE ) ),
	DefaultDelay=>VitalZeroDelay01,
	Mode=>VitalInertial,
	XON=>TRUE,
	MsgOn=>TRUE,
	MsgSeverity=>WARNING );

 VitalPathDelay01Z ( IO, IOGLITCH_DATA, "IO", IO_zd,
	Paths => (
	0 => ( OE_ipd'LAST_EVENT, tpd_OE_IO, TRUE ),
        1 => ( CLK_dly'LAST_EVENT, tpd_CLK_IO, TRUE ),
        2 => ( S_CLK_dly'LAST_EVENT, tpd_S_IO, TRUE ) ),
	DefaultDelay=>VitalZeroDelay01Z,
	Mode=>VitalInertial,
	XON=>TRUE,
	MsgOn=>TRUE,
	MsgSeverity=>WARNING );


END PROCESS VitalBehaviour_1;
END VITAL_VF;
configuration CFG_ROLIS_VITAL of ROLIS is 
        for VITAL_VF
        end for; 
end CFG_ROLIS_VITAL;
---------------------------------------------------------------------------------
-- VITAL model for cell RORI
---------------------------------------------------------------------------------
LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.VITAL_timing.all;
USE IEEE.VITAL_primitives.all;
LIBRARY VF1;
USE VF1.VLOGTOVITAL_TABLES.all;
-----------------------------------------------------------------------------
--ENTITY DECLARATION
-----------------------------------------------------------------------------
ENTITY RORI IS

GENERIC (
	tipd_IO			 : VITALDELAYTYPE01Z 	 := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
	tipd_D			 : VITALDELAYTYPE01Z 	 := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
	tipd_CLKI		 : VITALDELAYTYPE01Z 	 := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
	tipd_CLKO		 : VITALDELAYTYPE01Z 	 := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
	tipd_OE			 : VITALDELAYTYPE01Z 	 := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
	TimingChecksOn           : BOOLEAN               := TRUE;
	ticd_CLKO		 : VITALDELAYTYPE 	 := 0 ns;
	tisd_D_CLKO		 : VITALDELAYTYPE 	 := 0 ns;
	Xon                      : BOOLEAN               := TRUE;
	InstancePath             : STRING                := "*";
	MsgOn                    : BOOLEAN               := TRUE;
	tsetup_D_CLKO_noedge_posedge : VITALDELAYTYPE 	 := 0.36 ns;
	thold_D_CLKO_noedge_posedge : VITALDELAYTYPE 	 := 0.56 ns;
	tpw_CLKO_posedge : VITALDELAYTYPE 	 := 0.72 ns;
	tpw_CLKO_negedge : VITALDELAYTYPE 	 := 0 ns;
	tperiod_CLKO_posedge : VITALDELAYTYPE 	 := 1.44 ns;
	ticd_CLKI		 : VITALDELAYTYPE 	 := 0 ns;
	tpw_CLKI_posedge	 : VITALDELAYTYPE 	 := 0.66 ns;
	tpw_CLKI_negedge	 : VITALDELAYTYPE 	 := 0 ns;
	tperiod_CLKI_posedge	 : VITALDELAYTYPE 	 := 1.32 ns;
	tisd_IO_CLKI		 : VITALDELAYTYPE 	 := 0 ns;
	tsetup_IO_CLKI_noedge_posedge : VITALDELAYTYPE 	 := 0.33 ns;
	thold_IO_CLKI_noedge_posedge : VITALDELAYTYPE 	 := 0.53 ns;
	tpd_OE_IO		 : VITALDELAYTYPE01Z 	 := (0.64 ns, 0.64 ns, 0.64 ns, 0.64 ns, 0.64 ns, 0.64 ns);
	tpd_IO_O		 : VITALDELAYTYPE01 	 := (0.4 ns, 0.4 ns);
	tpd_CLKO_O		 : VITALDELAYTYPE01 	 := (3.14 ns, 3.14 ns);
	tpd_CLKO_IO		 : VITALDELAYTYPE01Z 	 := (2.74 ns, 2.74 ns, 2.74 ns, 2.74 ns, 2.74 ns, 2.74 ns);
	tpd_CLKI_Q		 : VITALDELAYTYPE01 	 := (1.23 ns, 1.23 ns)
	);

PORT    (
	O			 : OUT   std_logic;
	Q			 : OUT   std_logic;
	IO			 : INOUT std_logic := 'U';
	D			 : IN    std_logic := 'U';
	CLKI			 : IN    std_logic := 'U';
	CLKO			 : IN    std_logic := 'U';
	OE			 : IN    std_logic := 'U'
	);

ATTRIBUTE VITAL_LEVEL0 OF RORI : ENTITY IS TRUE ;

END RORI;

-----------------------------------------------------------------------------
-- ARCHITECTURE declaration
-----------------------------------------------------------------------------
ARCHITECTURE VITAL_VF OF RORI  IS
	ATTRIBUTE VITAL_LEVEL1 OF VITAL_VF : ARCHITECTURE IS TRUE;

	SIGNAL	IO_ipd			 : std_ulogic         := 'X';
	SIGNAL	D_ipd			 : std_ulogic         := 'X';
	SIGNAL	CLKI_ipd		 : std_ulogic         := 'X';
	SIGNAL	CLKO_ipd		 : std_ulogic         := 'X';
	SIGNAL	OE_ipd			 : std_ulogic         := 'X';
	SIGNAL	CLKI_dly		 : std_ulogic        := 'X';
	SIGNAL	D_dly			 : std_ulogic        := 'X';
	SIGNAL	CLKO_dly		 : std_ulogic        := 'X';
	SIGNAL	IO_dly			 : std_ulogic        := 'X';
BEGIN
-----------------------------------------------------------------------------
-- INPUT PATH DELAYs
-----------------------------------------------------------------------------
WIREDELAY : BLOCK
BEGIN
	VitalWireDelay( IO_ipd, IO, tipd_IO );
	VitalWireDelay( D_ipd, D, tipd_D );
	VitalWireDelay( CLKI_ipd, CLKI, tipd_CLKI );
	VitalWireDelay( CLKO_ipd, CLKO, tipd_CLKO );
	VitalWireDelay( OE_ipd, OE, tipd_OE );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
	VitalSignalDelay ( CLKI_dly, CLKI_ipd, ticd_CLKI);
	VitalSignalDelay ( D_dly, D_ipd, tisd_D_CLKO);
	VitalSignalDelay ( CLKO_dly, CLKO_ipd, ticd_CLKO);
	VitalSignalDelay ( IO_dly, IO_ipd, tisd_IO_CLKI);
END BLOCK;

-----------------------------------------------------------------------------
-- Behavior Section
-----------------------------------------------------------------------------

VitalBehaviour_0 : PROCESS(OE_ipd,D_dly,CLKO_dly,IO_dly,CLKI_dly)

VARIABLE 	Tviol_CLKO_D_flag1	 : std_ulogic		 := '0';
VARIABLE 	TimingData_D_CLKO1	 : VitalTimingDataType	 := VitalTimingDataInit;
VARIABLE 	Tviol_CLKO_flag2	 : std_ulogic		 := '0';
VARIABLE 	PeriodData_CLKO2	 : VitalPeriodDataType	 := VitalPeriodDataInit;
VARIABLE 	Tviol_CLKO_flag3	 : std_ulogic		 := '0';
VARIABLE 	PeriodData_CLKO3	 : VitalPeriodDataType	 := VitalPeriodDataInit;
VARIABLE 	Tviol_CLKI_flag4	 : std_ulogic		 := '0';
VARIABLE 	PeriodData_CLKI4	 : VitalPeriodDataType	 := VitalPeriodDataInit;
VARIABLE 	Tviol_CLKI_flag5	 : std_ulogic		 := '0';
VARIABLE 	PeriodData_CLKI5	 : VitalPeriodDataType	 := VitalPeriodDataInit;
VARIABLE 	Tviol_CLKI_IO_flag6	 : std_ulogic		 := '0';
VARIABLE 	TimingData_IO_CLKI6	 : VitalTimingDataType	 := VitalTimingDataInit;
VARIABLE 	Q_int_zd		 : std_ulogic;
VARIABLE 	VCC_zd			 : std_ulogic;
VARIABLE 	notifier_zd		 : std_ulogic;
VARIABLE 	PrevDataIn0		 : std_logic_vector (0 to 3) ;
VARIABLE 	Q_zd			 : std_ulogic;
VARIABLE 	PrevDataIn1		 : std_logic_vector (0 to 3) ;
VARIABLE 	IO_zd			 : std_ulogic;
VARIABLE 	O_zd			 : std_ulogic;
VARIABLE 	OGLITCH_DATA		 : VitalGlitchDataType;
VARIABLE 	QGLITCH_DATA		 : VitalGlitchDataType;
VARIABLE 	IOGLITCH_DATA		 : VitalGlitchDataType;
VARIABLE 	Violation_Flag		 : std_ulogic;


BEGIN

--Timing Check Section

IF(TimingChecksOn) THEN
VitalSetupHoldCheck(Violation => Tviol_CLKO_D_flag1,
TimingData => TimingData_D_CLKO1,
TestSignal => D_dly,
TestSignalName => "D",
TestDelay => 0 ns,
RefSignal => CLKO_dly,
RefSignalName => "CLKO",
RefDelay => 0 ns,
SetupHigh => tsetup_D_CLKO_noedge_posedge,
SetupLow => tsetup_D_CLKO_noedge_posedge,
HoldHigh => thold_D_CLKO_noedge_posedge,
HoldLow => thold_D_CLKO_noedge_posedge,
CheckEnabled => ( To_X01( OE_ipd )= '1' ),
RefTransition => '/',
HeaderMsg => InstancePath & "/RORI",
Xon => Xon,
MsgOn => MsgOn,
MsgSeverity => WARNING);


VitalPeriodPulseCheck(Violation => Tviol_CLKO_flag2,
PeriodData => PeriodData_CLKO2,
TestSignal => CLKO_dly,
TestSignalName => "CLKO",
TestDelay => 0 ns,
Period => 0 ns,
PulseWidthHigh => tpw_CLKO_posedge,
PulseWidthLow => tpw_CLKO_negedge,
CheckEnabled => ( To_X01( OE_ipd )= '1' ),
HeaderMsg => InstancePath & "/RORI",
Xon => Xon,
MsgOn => MsgOn,
MsgSeverity => WARNING);


VitalPeriodPulseCheck(Violation => Tviol_CLKO_flag3,
PeriodData => PeriodData_CLKO3,
TestSignal => CLKO_dly,
TestSignalName => "CLKO",
TestDelay => 0 ns,
Period => tperiod_CLKO_posedge,
PulseWidthHigh => 0 ns,
PulseWidthLow => 0 ns,
CheckEnabled => posedge( CLKO_dly'LAST_VALUE, CLKO_dly ) AND ( To_X01( OE_ipd )= '1' ),
HeaderMsg => InstancePath & "/RORI",
Xon => Xon,
MsgOn => MsgOn,
MsgSeverity => WARNING);


VitalPeriodPulseCheck(Violation => Tviol_CLKI_flag4,
PeriodData => PeriodData_CLKI4,
TestSignal => CLKI_dly,
TestSignalName => "CLKI",
TestDelay => 0 ns,
Period => 0 ns,
PulseWidthHigh => tpw_CLKI_posedge,
PulseWidthLow => tpw_CLKI_negedge,
CheckEnabled => TRUE,
HeaderMsg => InstancePath & "/RORI",
Xon => Xon,
MsgOn => MsgOn,
MsgSeverity => WARNING);


VitalPeriodPulseCheck(Violation => Tviol_CLKI_flag5,
PeriodData => PeriodData_CLKI5,
TestSignal => CLKI_dly,
TestSignalName => "CLKI",
TestDelay => 0 ns,
Period => tperiod_CLKI_posedge,
PulseWidthHigh => 0 ns,
PulseWidthLow => 0 ns,
CheckEnabled => posedge( CLKI_dly'LAST_VALUE, CLKI_dly ),
HeaderMsg => InstancePath & "/RORI",
Xon => Xon,
MsgOn => MsgOn,
MsgSeverity => WARNING);


VitalSetupHoldCheck(Violation => Tviol_CLKI_IO_flag6,
TimingData => TimingData_IO_CLKI6,
TestSignal => IO_dly,
TestSignalName => "IO",
TestDelay => 0 ns,
RefSignal => CLKI_dly,
RefSignalName => "CLKI",
RefDelay => 0 ns,
SetupHigh => tsetup_IO_CLKI_noedge_posedge,
SetupLow => tsetup_IO_CLKI_noedge_posedge,
HoldHigh => thold_IO_CLKI_noedge_posedge,
HoldLow => thold_IO_CLKI_noedge_posedge,
CheckEnabled => TRUE,
RefTransition => '/',
HeaderMsg => InstancePath & "/RORI",
Xon => Xon,
MsgOn => MsgOn,
MsgSeverity => WARNING);


END IF;   -- Timing Check Section

--Functionality Section

Violation_Flag	 := (((((Tviol_CLKO_D_flag1 or Tviol_CLKO_flag2) or Tviol_CLKO_flag3) or Tviol_CLKI_flag4) or Tviol_CLKI_flag5) or Tviol_CLKI_IO_flag6) ;
notifier_zd	 := 'X';
VitalStateTable(
StateTable => dfftab,
DataIn => std_logic_vector'(D_dly,CLKO_dly,'1','1'),
Result => Q_int_zd	,
PreviousDataIn => PrevDataIn0);

Q_int_zd	 := (Violation_Flag xor Q_int_zd);
IO_zd		 := VitalBUFIF1(Q_int_zd, OE_ipd);
O_zd		 := VitalBUF(IO_dly);
VitalStateTable(
StateTable => dfftab,
DataIn => std_logic_vector'(IO_dly,CLKI_dly,'1','1'),
Result => Q_zd		,
PreviousDataIn => PrevDataIn1);

Q_zd		 := (Violation_Flag xor Q_zd) ;

--PathDelay Section

 VitalPathDelay01 ( O, OGLITCH_DATA, "O", O_zd,
	Paths => (
	0 => ( IO_dly'LAST_EVENT, tpd_IO_O, TRUE ),
	1 => ( CLKO_dly'LAST_EVENT, tpd_CLKO_O, TRUE ) ),
	DefaultDelay=>VitalZeroDelay01,
	Mode=>VitalInertial,
	XON=>TRUE,
	MsgOn=>TRUE,
	MsgSeverity=>WARNING );

 VitalPathDelay01 ( Q, QGLITCH_DATA, "Q", Q_zd,
	Paths => (
	0 => ( CLKI_dly'LAST_EVENT, tpd_CLKI_Q, TRUE ) ),
	DefaultDelay=>VitalZeroDelay01,
	Mode=>VitalInertial,
	XON=>TRUE,
	MsgOn=>TRUE,
	MsgSeverity=>WARNING );

 VitalPathDelay01Z ( IO, IOGLITCH_DATA, "IO", IO_zd,
	Paths => (
	0 => ( OE_ipd'LAST_EVENT, VitalExtendToFillDelay(tpd_OE_IO), TRUE ),
	1 => ( CLKO_dly'LAST_EVENT, VitalExtendToFillDelay(tpd_CLKO_IO), TRUE ) ),
	DefaultDelay=>VitalZeroDelay01Z,
	Mode=>VitalInertial,
	XON=>TRUE,
	MsgOn=>TRUE,
	MsgSeverity=>WARNING );







END PROCESS VitalBehaviour_0;


END VITAL_VF;
configuration CFG_RORI_VITAL of RORI is 
        for VITAL_VF
        end for; 
end CFG_RORI_VITAL;
---------------------------------------------------------------------------------
-- VITAL model for cell RORIR
---------------------------------------------------------------------------------
LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.VITAL_timing.all;
USE IEEE.VITAL_primitives.all;
LIBRARY VF1;
USE VF1.all;
USE VF1.VLOGTOVITAL_TABLES.all;
-----------------------------------------------------------------------------
--ENTITY DECLARATION
-----------------------------------------------------------------------------
ENTITY RORIR IS

GENERIC (
	tipd_IO			 : VITALDELAYTYPE01Z 	 := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
	tipd_D			 : VITALDELAYTYPE01Z 	 := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
	tipd_CLKI		 : VITALDELAYTYPE01Z 	 := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
	tipd_CLKO		 : VITALDELAYTYPE01Z 	 := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
	tipd_OE			 : VITALDELAYTYPE01Z 	 := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
	tipd_R			 : VITALDELAYTYPE01Z 	 := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
	TimingChecksOn           : BOOLEAN               := TRUE;
	ticd_CLKO		 : VITALDELAYTYPE 	 := 0 ns;
	tisd_D_CLKO		 : VITALDELAYTYPE 	 := 0 ns;
	Xon                      : BOOLEAN               := TRUE;
	InstancePath             : STRING                := "*";
	MsgOn                    : BOOLEAN               := TRUE;
	tsetup_D_CLKO_noedge_posedge : VITALDELAYTYPE 	 := 0.36 ns;
	thold_D_CLKO_noedge_posedge : VITALDELAYTYPE 	 := 0.56 ns;
	tpw_CLKO_posedge : VITALDELAYTYPE 	 := 0.72 ns;
	tpw_CLKO_negedge : VITALDELAYTYPE 	 := 0 ns;
	tperiod_CLKO_posedge : VITALDELAYTYPE 	 := 1.44 ns;
	tisd_R_CLKO			 : VITALDELAYTYPE 	 := 0 ns;
	trecovery_CLKO_R_posedge_posedge : VITALDELAYTYPE 	 := 0.33 ns;
	tremoval_CLKO_R_posedge_posedge : VITALDELAYTYPE 	 := 0.53 ns;
	ticd_CLKI		 : VITALDELAYTYPE 	 := 0 ns;
	tisd_IO_CLKI		 : VITALDELAYTYPE 	 := 0 ns;
	tsetup_IO_CLKI_noedge_posedge : VITALDELAYTYPE 	 := 0.33 ns;
	thold_IO_CLKI_noedge_posedge : VITALDELAYTYPE 	 := 0.53 ns;
	tpw_CLKI_posedge	 : VITALDELAYTYPE 	 := 0.66 ns;
	tpw_CLKI_negedge	 : VITALDELAYTYPE 	 := 0 ns;
	tperiod_CLKI_posedge	 : VITALDELAYTYPE 	 := 1.32 ns;
	tisd_R_CLKI			 : VITALDELAYTYPE 	 := 0 ns;
	trecovery_CLKI_R_posedge_posedge : VITALDELAYTYPE 	 := 0.33 ns;
	tremoval_CLKI_R_posedge_posedge : VITALDELAYTYPE 	 := 0.53 ns;
	tpd_OE_IO		 : VITALDELAYTYPE01Z 	 := (0.64 ns, 0.64 ns, 0.64 ns, 0.64 ns, 0.64 ns, 0.64 ns);
	tpd_IO_O		 : VITALDELAYTYPE01 	 := (0.4 ns, 0.4 ns);
	tpd_CLKO_O		 : VITALDELAYTYPE01 	 := (3.14 ns, 3.14 ns);
	tpd_CLKO_IO		 : VITALDELAYTYPE01Z 	 := (2.74 ns, 2.74 ns, 2.74 ns, 2.74 ns, 2.74 ns, 2.74 ns);
	tpd_R_O			 : VITALDELAYTYPE01 	 := (3.14 ns, 3.14 ns);
	tbpd_R_O_CLKO			 : VITALDELAYTYPE01 	 := (3.14 ns, 3.14 ns);
	tpd_R_IO		 : VITALDELAYTYPE01Z 	 := (2.74 ns, 2.74 ns, 2.74 ns, 2.74 ns, 2.74 ns, 2.74 ns);
	tbpd_R_IO_CLKO		 : VITALDELAYTYPE01Z 	 := (2.74 ns, 2.74 ns, 2.74 ns, 2.74 ns, 2.74 ns, 2.74 ns);
	tpd_R_Q			 : VITALDELAYTYPE01 	 := (1.23 ns, 1.23 ns);
	tbpd_R_Q_CLKI			 : VITALDELAYTYPE01 	 := (1.23 ns, 1.23 ns);
	tpd_CLKI_Q		 : VITALDELAYTYPE01 	 := (1.23 ns, 1.23 ns)
	);

PORT    (
	O			 : OUT   std_logic;
	Q			 : OUT   std_logic;
	IO			 : INOUT std_logic := 'U';
	D			 : IN    std_logic := 'U';
	CLKI			 : IN    std_logic := 'U';
	CLKO			 : IN    std_logic := 'U';
	OE			 : IN    std_logic := 'U';
	R			 : IN    std_logic := 'U'
	);

ATTRIBUTE VITAL_LEVEL0 OF RORIR : ENTITY IS TRUE ;

END RORIR;

-----------------------------------------------------------------------------
-- ARCHITECTURE declaration
-----------------------------------------------------------------------------
ARCHITECTURE VITAL_VF OF RORIR  IS
	ATTRIBUTE VITAL_LEVEL1 OF VITAL_VF : ARCHITECTURE IS TRUE;

	SIGNAL	IO_ipd			 : std_logic         := 'X';
	SIGNAL	D_ipd			 : std_logic         := 'X';
	SIGNAL	CLKI_ipd		 : std_logic         := 'X';
	SIGNAL	CLKO_ipd		 : std_logic         := 'X';
	SIGNAL	OE_ipd			 : std_logic         := 'X';
	SIGNAL	R_ipd			 : std_logic         := 'X';
	SIGNAL	CLKI_dly		 : std_ulogic        := 'X';
	SIGNAL	D_dly			 : std_ulogic        := 'X';
	SIGNAL	R1_dly			 : std_ulogic        := 'X';
	SIGNAL	R2_dly			 : std_ulogic        := 'X';
	SIGNAL	CLKO_dly		 : std_ulogic        := 'X';
	SIGNAL	IO_dly			 : std_ulogic        := 'X';
BEGIN
-----------------------------------------------------------------------------
-- INPUT PATH DELAYs
-----------------------------------------------------------------------------
WIREDELAY : BLOCK
BEGIN
	VitalWireDelay( IO_ipd, IO, tipd_IO );
	VitalWireDelay( D_ipd, D, tipd_D );
	VitalWireDelay( CLKI_ipd, CLKI, tipd_CLKI );
	VitalWireDelay( CLKO_ipd, CLKO, tipd_CLKO );
	VitalWireDelay( OE_ipd, OE, tipd_OE );
	VitalWireDelay( R_ipd, R, tipd_R );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
	VitalSignalDelay ( CLKI_dly, CLKI_ipd, ticd_CLKI);
	VitalSignalDelay ( D_dly, D_ipd, tisd_D_CLKO);
	VitalSignalDelay ( R1_dly, R_ipd, tisd_R_CLKO);
	VitalSignalDelay ( R2_dly, R_ipd, tisd_R_CLKi);
	VitalSignalDelay ( CLKO_dly, CLKO_ipd, ticd_CLKO);
	VitalSignalDelay ( IO_dly, IO_ipd, tisd_IO_CLKI);
END BLOCK;

-----------------------------------------------------------------------------
-- Behavior Section
-----------------------------------------------------------------------------

VitalBehaviour_0 : PROCESS(OE_ipd,D_dly,CLKO_dly,R1_dly,R2_dly,IO_dly,CLKI_dly)

VARIABLE 	Tviol_CLKO_D_flag1	 : std_ulogic		 := '0';
VARIABLE 	TimingData_D_CLKO1	 : VitalTimingDataType	 := VitalTimingDataInit;
VARIABLE 	Tviol_CLKO_flag2	 : std_ulogic		 := '0';
VARIABLE 	PeriodData_CLKO2	 : VitalPeriodDataType	 := VitalPeriodDataInit;
VARIABLE 	Tviol_CLKO_flag3	 : std_ulogic		 := '0';
VARIABLE 	PeriodData_CLKO3	 : VitalPeriodDataType	 := VitalPeriodDataInit;
VARIABLE 	Tviol_R_CLKO_flag4	 : std_ulogic		 := '0';
VARIABLE 	TimingData_CLKO_R4	 : VitalTimingDataType	 := VitalTimingDataInit;
VARIABLE 	Tviol_R_CLKI_flag4	 : std_ulogic		 := '0';
VARIABLE 	TimingData_CLKI_R4	 : VitalTimingDataType	 := VitalTimingDataInit;
VARIABLE 	Tviol_CLKI_IO_flag6	 : std_ulogic		 := '0';
VARIABLE 	TimingData_IO_CLKI6	 : VitalTimingDataType	 := VitalTimingDataInit;
VARIABLE 	Tviol_CLKI_flag7	 : std_ulogic		 := '0';
VARIABLE 	PeriodData_CLKI7	 : VitalPeriodDataType	 := VitalPeriodDataInit;
VARIABLE 	Tviol_CLKI_flag8	 : std_ulogic		 := '0';
VARIABLE 	PeriodData_CLKI8	 : VitalPeriodDataType	 := VitalPeriodDataInit;
VARIABLE 	Q_int_zd		 : std_ulogic;
VARIABLE 	VCC_zd			 : std_ulogic;
VARIABLE 	Bool_SenseList		 : BOOLEAN;
VARIABLE 	notifier_zd		 : std_ulogic;
VARIABLE 	PrevDataIn0		 : std_logic_vector (0 to 3) ;
VARIABLE 	Q_zd			 : std_ulogic;
VARIABLE 	PrevDataIn1		 : std_logic_vector (0 to 3) ;
VARIABLE 	OE_R_zd		 : std_ulogic;
VARIABLE 	IO_zd			 : std_ulogic;
VARIABLE 	O_zd			 : std_ulogic;
VARIABLE 	OGLITCH_DATA		 : VitalGlitchDataType;
VARIABLE 	QGLITCH_DATA		 : VitalGlitchDataType;
VARIABLE 	IOGLITCH_DATA		 : VitalGlitchDataType;
VARIABLE 	Violation_Flag		 : std_ulogic;


BEGIN

--Timing Check Section

IF(TimingChecksOn) THEN
VitalSetupHoldCheck(Violation => Tviol_CLKO_D_flag1,
TimingData => TimingData_D_CLKO1,
TestSignal => D_dly,
TestSignalName => "D",
TestDelay => 0 ns,
RefSignal => CLKO_dly,
RefSignalName => "CLKO",
RefDelay => 0 ns,
SetupHigh => tsetup_D_CLKO_noedge_posedge,
SetupLow => tsetup_D_CLKO_noedge_posedge,
HoldHigh => thold_D_CLKO_noedge_posedge,
HoldLow => thold_D_CLKO_noedge_posedge,
CheckEnabled => ( To_X01( OE_R_zd )= '1' ),
RefTransition => '/',
HeaderMsg => InstancePath & "/RORIR",
Xon => Xon,
MsgOn => MsgOn,
MsgSeverity => WARNING);


VitalPeriodPulseCheck(Violation => Tviol_CLKO_flag2,
PeriodData => PeriodData_CLKO2,
TestSignal => CLKO_dly,
TestSignalName => "CLKO",
TestDelay => 0 ns,
Period => 0 ns,
PulseWidthHigh => tpw_CLKO_posedge,
PulseWidthLow => tpw_CLKO_negedge,
CheckEnabled => ( To_X01( OE_R_zd )= '1' ),
HeaderMsg => InstancePath & "/RORIR",
Xon => Xon,
MsgOn => MsgOn,
MsgSeverity => WARNING);


VitalPeriodPulseCheck(Violation => Tviol_CLKO_flag3,
PeriodData => PeriodData_CLKO3,
TestSignal => CLKO_dly,
TestSignalName => "CLKO",
TestDelay => 0 ns,
Period => tperiod_CLKO_posedge,
PulseWidthHigh => 0 ns,
PulseWidthLow => 0 ns,
CheckEnabled => posedge( CLKO_dly'LAST_VALUE, CLKO_dly ) AND ( To_X01( OE_R_zd )= '1' ),
HeaderMsg => InstancePath & "/RORIR",
Xon => Xon,
MsgOn => MsgOn,
MsgSeverity => WARNING);


VitalRecoveryRemovalCheck(Violation => Tviol_R_CLKO_flag4,
TimingData => TimingData_CLKO_R4,
TestSignal => CLKO_dly,
TestSignalName => "CLKO",
TestDelay => 0 ns,
RefSignal => R1_dly,
RefSignalName => "R",
RefDelay => 0 ns,
Recovery => trecovery_CLKO_R_posedge_posedge,
Removal => tremoval_CLKO_R_posedge_posedge,
ActiveLow => FALSE,
CheckEnabled => ( To_X01( OE_ipd )= '1' ),
RefTransition => '/',
HeaderMsg =>InstancePath & "/RORIR",
Xon => Xon,
MsgOn => MsgOn,
MsgSeverity => WARNING);




VitalSetupHoldCheck(Violation => Tviol_CLKI_IO_flag6,
TimingData => TimingData_IO_CLKI6,
TestSignal => IO_dly,
TestSignalName => "IO",
TestDelay => 0 ns,
RefSignal => CLKI_dly,
RefSignalName => "CLKI",
RefDelay => 0 ns,
SetupHigh => tsetup_IO_CLKI_noedge_posedge,
SetupLow => tsetup_IO_CLKI_noedge_posedge,
HoldHigh => thold_IO_CLKI_noedge_posedge,
HoldLow => thold_IO_CLKI_noedge_posedge,
CheckEnabled => ( To_X01( R2_dly )= '0' ),
RefTransition => '/',
HeaderMsg => InstancePath & "/RORIR",
Xon => Xon,
MsgOn => MsgOn,
MsgSeverity => WARNING);


VitalPeriodPulseCheck(Violation => Tviol_CLKI_flag7,
PeriodData => PeriodData_CLKI7,
TestSignal => CLKI_dly,
TestSignalName => "CLKI",
TestDelay => 0 ns,
Period => 0 ns,
PulseWidthHigh => tpw_CLKI_posedge,
PulseWidthLow => tpw_CLKI_negedge,
CheckEnabled => ( To_X01( R2_dly )= '0' ),
HeaderMsg => InstancePath & "/RORIR",
Xon => Xon,
MsgOn => MsgOn,
MsgSeverity => WARNING);


VitalPeriodPulseCheck(Violation => Tviol_CLKI_flag8,
PeriodData => PeriodData_CLKI8,
TestSignal => CLKI_dly,
TestSignalName => "CLKI",
TestDelay => 0 ns,
Period => tperiod_CLKI_posedge,
PulseWidthHigh => 0 ns,
PulseWidthLow => 0 ns,
CheckEnabled => posedge( CLKI_dly'LAST_VALUE, CLKI_dly ) AND ( To_X01( R2_dly )= '0' ),
HeaderMsg => InstancePath & "/RORIR",
Xon => Xon,
MsgOn => MsgOn,
MsgSeverity => WARNING);

VitalRecoveryRemovalCheck(Violation => Tviol_R_CLKI_flag4,
TimingData => TimingData_CLKI_R4,
TestSignal => CLKI_dly,
TestSignalName => "CLKI",
TestDelay => 0 ns,
RefSignal => R2_dly,
RefSignalName => "R",
RefDelay => 0 ns,
Recovery => trecovery_CLKI_R_posedge_posedge,
Removal => tremoval_CLKI_R_posedge_posedge,
ActiveLow => FALSE,
CheckEnabled => TRUE,
RefTransition => '/',
HeaderMsg =>InstancePath & "/RORIR",
Xon => Xon,
MsgOn => MsgOn,
MsgSeverity => WARNING);


END IF;   -- Timing Check Section

--Functionality Section

Violation_Flag	 := ((((((Tviol_CLKO_D_flag1 or Tviol_CLKO_flag2)
 or Tviol_CLKO_flag3)
 or Tviol_R_CLKO_flag4
 or Tviol_R_CLKI_flag4)
 or Tviol_CLKI_IO_flag6)
 or Tviol_CLKI_flag7)
 or Tviol_CLKI_flag8)
;
VCC_zd		 := '1';
notifier_zd	 := 'X';
VitalStateTable(
StateTable => dfftab,
DataIn => std_logic_vector'(D_dly,CLKO_dly,NOT(R1_dly),VCC_zd),
Result => Q_int_zd	,
PreviousDataIn => PrevDataIn0);

Q_int_zd	 := (Violation_Flag xor Q_int_zd);
IO_zd		 := VitalBUFIF1(Q_int_zd,OE_ipd);


O_zd		 := VitalBUF(IO_dly);

VitalStateTable(
StateTable => dfftab,
DataIn => std_logic_vector'(IO_dly,CLKI_dly,NOT(R2_dly),VCC_zd),
Result => Q_zd		,
PreviousDataIn => PrevDataIn1);

OE_R_zd	 := VitalAND2(OE_ipd,NOT(R1_dly));
Q_zd		 := (Violation_Flag xor Q_zd);

--PathDelay Section

 VitalPathDelay01 ( O, OGLITCH_DATA, "O", O_zd,
	Paths => (
	0 => ( IO_dly'LAST_EVENT, tpd_IO_O, TRUE ),
	1 => ( CLKO_dly'LAST_EVENT, tpd_CLKO_O, TRUE ),
	2 => ( R1_dly'LAST_EVENT, tbpd_R_O_CLKO, TRUE ) ),
	DefaultDelay=>VitalZeroDelay01,
	Mode=>VitalInertial,
	XON=>TRUE,
	MsgOn=>TRUE,
	MsgSeverity=>WARNING );

 VitalPathDelay01 ( Q, QGLITCH_DATA, "Q", Q_zd,
	Paths => (
	0 => ( CLKI_dly'LAST_EVENT, tpd_CLKI_Q, TRUE ),
        1 => ( R2_dly'LAST_EVENT, tbpd_R_Q_CLKI, TRUE ) ),
	DefaultDelay=>VitalZeroDelay01,
	Mode=>VitalInertial,
	XON=>TRUE,
	MsgOn=>TRUE,
	MsgSeverity=>WARNING );

 VitalPathDelay01Z ( IO, IOGLITCH_DATA, "IO", IO_zd,
	Paths => (
	0 => ( OE_ipd'LAST_EVENT, VitalExtendToFillDelay(tpd_OE_IO), TRUE ),
	1 => ( CLKO_dly'LAST_EVENT, VitalExtendToFillDelay(tpd_CLKO_IO), TRUE ),
	2 => ( R1_dly'LAST_EVENT, VitalExtendToFillDelay(tbpd_R_IO_CLKO), TRUE ) ),
	DefaultDelay=>VitalZeroDelay01Z,
	Mode=>VitalInertial,
	XON=>TRUE,
	MsgOn=>TRUE,
	MsgSeverity=>WARNING );




END PROCESS VitalBehaviour_0;


END VITAL_VF;
configuration CFG_RORIR_VITAL of RORIR is 
        for VITAL_VF
        end for; 
end CFG_RORIR_VITAL;
---------------------------------------------------------------------------------
-- VITAL model for cell RORIS
---------------------------------------------------------------------------------
LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.VITAL_timing.all;
USE IEEE.VITAL_primitives.all;
LIBRARY VF1;
USE VF1.all;
USE VF1.VLOGTOVITAL_TABLES.all;
-----------------------------------------------------------------------------
--ENTITY DECLARATION
-----------------------------------------------------------------------------
ENTITY RORIS IS

GENERIC (
	tipd_IO			 : VITALDELAYTYPE01Z 	 := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
	tipd_D			 : VITALDELAYTYPE01Z 	 := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
	tipd_CLKI		 : VITALDELAYTYPE01Z 	 := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
	tipd_CLKO		 : VITALDELAYTYPE01Z 	 := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
	tipd_OE			 : VITALDELAYTYPE01Z 	 := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
	tipd_S			 : VITALDELAYTYPE01Z 	 := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
	TimingChecksOn           : BOOLEAN               := TRUE;
	ticd_CLKO		 : VITALDELAYTYPE 	 := 0 ns;
	tisd_D_CLKO		 : VITALDELAYTYPE 	 := 0 ns;
	Xon                      : BOOLEAN               := TRUE;
	InstancePath             : STRING                := "*";
	MsgOn                    : BOOLEAN               := TRUE;
	tsetup_D_CLKO_noedge_posedge : VITALDELAYTYPE 	 := 0.36 ns;
	thold_D_CLKO_noedge_posedge : VITALDELAYTYPE 	 := 0.56 ns;
	tpw_CLKO_posedge : VITALDELAYTYPE 	 := 0.72 ns;
	tpw_CLKO_negedge : VITALDELAYTYPE 	 := 0 ns;
	tperiod_CLKO_posedge : VITALDELAYTYPE 	 := 1.44 ns;
	tisd_S_CLKO			 : VITALDELAYTYPE 	 := 0 ns;
	trecovery_CLKO_S_posedge_posedge : VITALDELAYTYPE 	 := 0.33 ns;
	tremoval_CLKO_S_posedge_posedge : VITALDELAYTYPE 	 := 0.53 ns;
	ticd_CLKI		 : VITALDELAYTYPE 	 := 0 ns;
	tisd_IO_CLKI		 : VITALDELAYTYPE 	 := 0 ns;
	tsetup_IO_CLKI_noedge_posedge : VITALDELAYTYPE 	 := 0.33 ns;
	thold_IO_CLKI_noedge_posedge : VITALDELAYTYPE 	 := 0.53 ns;
	tpw_CLKI_posedge	 : VITALDELAYTYPE 	 := 0.66 ns;
	tpw_CLKI_negedge	 : VITALDELAYTYPE 	 := 0 ns;
	tperiod_CLKI_posedge	 : VITALDELAYTYPE 	 := 1.32 ns;
	tisd_S_CLKI			 : VITALDELAYTYPE 	 := 0 ns;
	trecovery_CLKI_S_posedge_posedge : VITALDELAYTYPE 	 := 0.33 ns;
	tremoval_CLKI_S_posedge_posedge : VITALDELAYTYPE 	 := 0.53 ns;
	tpd_OE_IO		 : VITALDELAYTYPE01Z 	 := (0.64 ns, 0.64 ns, 0.64 ns, 0.64 ns, 0.64 ns, 0.64 ns);
	tpd_IO_O		 : VITALDELAYTYPE01 	 := (0.4 ns, 0.4 ns);
	tpd_CLKO_O		 : VITALDELAYTYPE01 	 := (3.14 ns, 3.14 ns);
	tpd_CLKO_IO		 : VITALDELAYTYPE01Z 	 := (2.74 ns, 2.74 ns, 2.74 ns, 2.74 ns, 2.74 ns, 2.74 ns);
	tpd_S_O			 : VITALDELAYTYPE01 	 := (3.14 ns, 3.14 ns);
	tbpd_S_O_CLKO			 : VITALDELAYTYPE01 	 := (3.14 ns, 3.14 ns);
	tpd_S_IO		 : VITALDELAYTYPE01Z 	 := (2.74 ns, 2.74 ns, 2.74 ns, 2.74 ns, 2.74 ns, 2.74 ns);
	tbpd_S_IO_CLKO		 : VITALDELAYTYPE01Z 	 := (2.74 ns, 2.74 ns, 2.74 ns, 2.74 ns, 2.74 ns, 2.74 ns);
	tpd_S_Q		         : VITALDELAYTYPE01 	 := (1.23 ns, 1.23 ns);
	tbpd_S_Q_CLKI		         : VITALDELAYTYPE01 	 := (1.23 ns, 1.23 ns);
	tpd_CLKI_Q		 : VITALDELAYTYPE01 	 := (1.23 ns, 1.23 ns)
	);

PORT    (
	O			 : OUT   std_logic;
	Q			 : OUT   std_logic;
	IO			 : INOUT std_logic := 'U';
	D			 : IN    std_logic := 'U';
	CLKI			 : IN    std_logic := 'U';
	CLKO			 : IN    std_logic := 'U';
	OE			 : IN    std_logic := 'U';
	S			 : IN    std_logic := 'U'
	);

ATTRIBUTE VITAL_LEVEL0 OF RORIS : ENTITY IS TRUE ;

END RORIS;

-----------------------------------------------------------------------------
-- ARCHITECTURE declaration
-----------------------------------------------------------------------------
ARCHITECTURE VITAL_VF OF RORIS  IS
	ATTRIBUTE VITAL_LEVEL1 OF VITAL_VF : ARCHITECTURE IS TRUE;

	SIGNAL	IO_ipd			 : std_logic         := 'X';
	SIGNAL	D_ipd			 : std_logic         := 'X';
	SIGNAL	CLKI_ipd		 : std_logic         := 'X';
	SIGNAL	CLKO_ipd		 : std_logic         := 'X';
	SIGNAL	OE_ipd			 : std_logic         := 'X';
	SIGNAL	S_ipd			 : std_logic         := 'X';
	SIGNAL	CLKI_dly		 : std_ulogic        := 'X';
	SIGNAL	D_dly			 : std_ulogic        := 'X';
	SIGNAL	S1_dly			 : std_ulogic        := 'X';
	SIGNAL	S2_dly			 : std_ulogic        := 'X';
	SIGNAL	CLKO_dly		 : std_ulogic        := 'X';
	SIGNAL	IO_dly			 : std_ulogic        := 'X';
BEGIN
-----------------------------------------------------------------------------
-- INPUT PATH DELAYs
-----------------------------------------------------------------------------
WIREDELAY : BLOCK
BEGIN
	VitalWireDelay( IO_ipd, IO, tipd_IO );
	VitalWireDelay( D_ipd, D, tipd_D );
	VitalWireDelay( CLKI_ipd, CLKI, tipd_CLKI );
	VitalWireDelay( CLKO_ipd, CLKO, tipd_CLKO );
	VitalWireDelay( OE_ipd, OE, tipd_OE );
	VitalWireDelay( S_ipd, S, tipd_S );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
	VitalSignalDelay ( CLKI_dly, CLKI_ipd, ticd_CLKI);
	VitalSignalDelay ( D_dly, D_ipd, tisd_D_CLKO);
	VitalSignalDelay ( S1_dly, S_ipd, tisd_S_CLKO);
	VitalSignalDelay ( S2_dly, S_ipd, tisd_S_CLKI);
	VitalSignalDelay ( CLKO_dly, CLKO_ipd, ticd_CLKO);
	VitalSignalDelay ( IO_dly, IO_ipd, tisd_IO_CLKI);
END BLOCK;

-----------------------------------------------------------------------------
-- Behavior Section
-----------------------------------------------------------------------------

VitalBehaviour_0 : PROCESS(OE_ipd,D_dly,CLKI_dly,S1_dly,S2_dly,IO_dly,CLKO_dly)

VARIABLE 	Tviol_CLKO_D_flag1	 : std_ulogic		 := '0';
VARIABLE 	TimingData_D_CLKO1	 : VitalTimingDataType	 := VitalTimingDataInit;
VARIABLE 	Tviol_CLKO_flag2	 : std_ulogic		 := '0';
VARIABLE 	PeriodData_CLKO2	 : VitalPeriodDataType	 := VitalPeriodDataInit;
VARIABLE 	Tviol_CLKO_flag3	 : std_ulogic		 := '0';
VARIABLE 	PeriodData_CLKO3	 : VitalPeriodDataType	 := VitalPeriodDataInit;
VARIABLE 	Tviol_S_CLKO_flag4	 : std_ulogic		 := '0';
VARIABLE 	TimingData_CLKO_S4	 : VitalTimingDataType	 := VitalTimingDataInit;
VARIABLE 	Tviol_S_CLKI_flag4	 : std_ulogic		 := '0';
VARIABLE 	TimingData_CLKI_S4	 : VitalTimingDataType	 := VitalTimingDataInit;
VARIABLE 	Tviol_CLKI_IO_flag6	 : std_ulogic		 := '0';
VARIABLE 	TimingData_IO_CLKI6	 : VitalTimingDataType	 := VitalTimingDataInit;
VARIABLE 	Tviol_CLKI_flag7	 : std_ulogic		 := '0';
VARIABLE 	PeriodData_CLKI7	 : VitalPeriodDataType	 := VitalPeriodDataInit;
VARIABLE 	Tviol_CLKI_flag8	 : std_ulogic		 := '0';
VARIABLE 	PeriodData_CLKI8	 : VitalPeriodDataType	 := VitalPeriodDataInit;
VARIABLE 	Q_int_zd		 : std_ulogic;
VARIABLE 	VCC_zd			 : std_ulogic;
VARIABLE 	Bool_SenseList		 : BOOLEAN;
VARIABLE 	notifier_zd		 : std_ulogic;
VARIABLE 	PrevDataIn0		 : std_logic_vector (0 to 3) ;
VARIABLE 	Q_zd			 : std_ulogic;
VARIABLE 	PrevDataIn1		 : std_logic_vector (0 to 3) ;
VARIABLE 	OE_S_zd		 : std_ulogic;
VARIABLE 	IO_zd			 : std_ulogic;
VARIABLE 	O_zd			 : std_ulogic;
VARIABLE 	OGLITCH_DATA		 : VitalGlitchDataType;
VARIABLE 	QGLITCH_DATA		 : VitalGlitchDataType;
VARIABLE 	IOGLITCH_DATA		 : VitalGlitchDataType;
VARIABLE 	Violation_Flag		 : std_ulogic;


BEGIN

--Timing Check Section

IF(TimingChecksOn) THEN
VitalSetupHoldCheck(Violation => Tviol_CLKO_D_flag1,
TimingData => TimingData_D_CLKO1,
TestSignal => D_dly,
TestSignalName => "D",
TestDelay => 0 ns,
RefSignal => CLKO_dly,
RefSignalName => "CLKO",
RefDelay => 0 ns,
SetupHigh => tsetup_D_CLKO_noedge_posedge,
SetupLow => tsetup_D_CLKO_noedge_posedge,
HoldHigh => thold_D_CLKO_noedge_posedge,
HoldLow => thold_D_CLKO_noedge_posedge,
CheckEnabled => ( To_X01( OE_S_zd )= '1' ),
RefTransition => '/',
HeaderMsg => InstancePath & "/RORIS",
Xon => Xon,
MsgOn => MsgOn,
MsgSeverity => WARNING);


VitalPeriodPulseCheck(Violation => Tviol_CLKO_flag2,
PeriodData => PeriodData_CLKO2,
TestSignal => CLKO_dly,
TestSignalName => "CLKO",
TestDelay => 0 ns,
Period => 0 ns,
PulseWidthHigh => tpw_CLKO_posedge,
PulseWidthLow => tpw_CLKO_negedge,
CheckEnabled => ( To_X01( OE_S_zd )= '1' ),
HeaderMsg => InstancePath & "/RORIS",
Xon => Xon,
MsgOn => MsgOn,
MsgSeverity => WARNING);


VitalPeriodPulseCheck(Violation => Tviol_CLKO_flag3,
PeriodData => PeriodData_CLKO3,
TestSignal => CLKO_dly,
TestSignalName => "CLKO",
TestDelay => 0 ns,
Period => tperiod_CLKO_posedge,
PulseWidthHigh => 0 ns,
PulseWidthLow => 0 ns,
CheckEnabled => posedge( CLKO_dly'LAST_VALUE, CLKO_dly ) AND ( To_X01( OE_S_zd )= '1' ),
HeaderMsg => InstancePath & "/RORIS",
Xon => Xon,
MsgOn => MsgOn,
MsgSeverity => WARNING);


VitalRecoveryRemovalCheck(Violation => Tviol_S_CLKO_flag4,
TimingData => TimingData_CLKO_S4,
TestSignal => CLKO_dly,
TestSignalName => "CLKO",
TestDelay => 0 ns,
RefSignal => S1_dly,
RefSignalName => "S",
RefDelay => 0 ns,
Recovery => trecovery_CLKO_S_posedge_posedge,
Removal => tremoval_CLKO_S_posedge_posedge,
ActiveLow => FALSE,
CheckEnabled => ( To_X01( OE_ipd )= '1' ),
RefTransition => '/',
HeaderMsg =>InstancePath & "/RORIS",
Xon => Xon,
MsgOn => MsgOn,
MsgSeverity => WARNING);




VitalSetupHoldCheck(Violation => Tviol_CLKI_IO_flag6,
TimingData => TimingData_IO_CLKI6,
TestSignal => IO_dly,
TestSignalName => "IO",
TestDelay => 0 ns,
RefSignal => CLKI_dly,
RefSignalName => "CLKI",
RefDelay => 0 ns,
SetupHigh => tsetup_IO_CLKI_noedge_posedge,
SetupLow => tsetup_IO_CLKI_noedge_posedge,
HoldHigh => thold_IO_CLKI_noedge_posedge,
HoldLow => thold_IO_CLKI_noedge_posedge,
CheckEnabled => ( To_X01( S2_dly )= '0' ),
RefTransition => '/',
HeaderMsg => InstancePath & "/RORIS",
Xon => Xon,
MsgOn => MsgOn,
MsgSeverity => WARNING);


VitalPeriodPulseCheck(Violation => Tviol_CLKI_flag7,
PeriodData => PeriodData_CLKI7,
TestSignal => CLKI_dly,
TestSignalName => "CLKI",
TestDelay => 0 ns,
Period => 0 ns,
PulseWidthHigh => tpw_CLKI_posedge,
PulseWidthLow => tpw_CLKI_negedge,
CheckEnabled => ( To_X01( S2_dly )= '0' ),
HeaderMsg => InstancePath & "/RORIS",
Xon => Xon,
MsgOn => MsgOn,
MsgSeverity => WARNING);


VitalPeriodPulseCheck(Violation => Tviol_CLKI_flag8,
PeriodData => PeriodData_CLKI8,
TestSignal => CLKI_dly,
TestSignalName => "CLKI",
TestDelay => 0 ns,
Period => tperiod_CLKI_posedge,
PulseWidthHigh => 0 ns,
PulseWidthLow => 0 ns,
CheckEnabled => posedge( CLKI_dly'LAST_VALUE, CLKI_dly ) AND ( To_X01( S2_dly )= '0' ),
HeaderMsg => InstancePath & "/RORIS",
Xon => Xon,
MsgOn => MsgOn,
MsgSeverity => WARNING);

VitalRecoveryRemovalCheck(Violation => Tviol_S_CLKI_flag4,
TimingData => TimingData_CLKI_S4,
TestSignal => CLKI_dly,
TestSignalName => "CLKI",
TestDelay => 0 ns,
RefSignal => S2_dly,
RefSignalName => "S",
RefDelay => 0 ns,
Recovery => trecovery_CLKI_S_posedge_posedge,
Removal => tremoval_CLKI_S_posedge_posedge,
ActiveLow => FALSE,
CheckEnabled => TRUE,
RefTransition => '/',
HeaderMsg =>InstancePath & "/RORIS",
Xon => Xon,
MsgOn => MsgOn,
MsgSeverity => WARNING);


END IF;   -- Timing Check Section

--Functionality Section

Violation_Flag	 := ((((((Tviol_CLKO_D_flag1 or Tviol_CLKO_flag2)
 or Tviol_CLKO_flag3)
 or Tviol_S_CLKO_flag4
 or Tviol_S_CLKI_flag4)
 or Tviol_CLKI_IO_flag6)
 or Tviol_CLKI_flag7)
 or Tviol_CLKI_flag8)
;
VCC_zd		 := '1';
notifier_zd	 := 'X';
VitalStateTable(
StateTable => dfftab,
DataIn => std_logic_vector'(D_dly,CLKO_dly,VCC_zd,NOT(S1_dly)),
Result => Q_int_zd	,
PreviousDataIn => PrevDataIn0);

Q_int_zd	 := (Violation_Flag xor Q_int_zd);
IO_zd		 := VitalBUFIF1(Q_int_zd,OE_ipd);
O_zd		 := VitalBUF(IO_dly);

VitalStateTable(
StateTable => dfftab,
DataIn => std_logic_vector'(IO_dly,CLKI_dly,VCC_zd,NOT(S2_dly)),
Result => Q_zd		,
PreviousDataIn => PrevDataIn1);

OE_S_zd	 := VitalAND2(OE_ipd,NOT(S1_dly));
Q_zd		 := (Violation_Flag xor Q_zd);

--PathDelay Section

 VitalPathDelay01 ( O, OGLITCH_DATA, "O", O_zd,
	Paths => (
	0 => ( IO_dly'LAST_EVENT, tpd_IO_O, TRUE ),
	1 => ( CLKO_dly'LAST_EVENT, tpd_CLKO_O, TRUE ),
	2 => ( S1_dly'LAST_EVENT, tbpd_S_O_CLKO, TRUE ) ),
	DefaultDelay=>VitalZeroDelay01,
	Mode=>VitalInertial,
	XON=>TRUE,
	MsgOn=>TRUE,
	MsgSeverity=>WARNING );

 VitalPathDelay01 ( Q, QGLITCH_DATA, "Q", Q_zd,
	Paths => (
	0 => ( CLKI_dly'LAST_EVENT, tpd_CLKI_Q, TRUE ),
        1 => ( S2_dly'LAST_EVENT, tbpd_S_Q_CLKI, TRUE ) ),
	DefaultDelay=>VitalZeroDelay01,
	Mode=>VitalInertial,
	XON=>TRUE,
	MsgOn=>TRUE,
	MsgSeverity=>WARNING );

 VitalPathDelay01Z ( IO, IOGLITCH_DATA, "IO", IO_zd,
	Paths => (
	0 => ( OE_ipd'LAST_EVENT, tpd_OE_IO, TRUE ),
	1 => ( CLKO_dly'LAST_EVENT, tpd_CLKO_IO, TRUE ),
	2 => ( S1_dly'LAST_EVENT, tbpd_S_IO_CLKO, TRUE ) ),
	DefaultDelay=>VitalZeroDelay01Z,
	Mode=>VitalInertial,
	XON=>TRUE,
	MsgOn=>TRUE,
	MsgSeverity=>WARNING );


END PROCESS VitalBehaviour_0;


END VITAL_VF;
configuration CFG_RORIS_VITAL of RORIS is 
        for VITAL_VF
        end for; 
end CFG_RORIS_VITAL;
---------------------------------------------------------------------------------
-- VITAL model for cell ROT
---------------------------------------------------------------------------------
LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.VITAL_timing.all;
USE IEEE.VITAL_primitives.all;
LIBRARY VF1;
USE VF1.VLOGTOVITAL_TABLES.all;
-----------------------------------------------------------------------------
--ENTITY DECLARATION
-----------------------------------------------------------------------------
ENTITY ROT IS

GENERIC (
	tipd_D			 : VITALDELAYTYPE01Z 	 := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
	tipd_CLK		 : VITALDELAYTYPE01Z 	 := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
	tipd_OE			 : VITALDELAYTYPE01Z 	 := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
	TimingChecksOn           : BOOLEAN               := TRUE;
	ticd_CLK		 : VITALDELAYTYPE 	 := 0 ns;
	tisd_D_CLK		 : VITALDELAYTYPE 	 := 0 ns;
	Xon                      : BOOLEAN               := TRUE;
	InstancePath             : STRING                := "*";
	MsgOn                    : BOOLEAN               := TRUE;
	tsetup_D_CLK_noedge_posedge : VITALDELAYTYPE 	 := 0.36 ns;
	thold_D_CLK_noedge_posedge : VITALDELAYTYPE 	 := 0.56 ns;
	tpw_CLK_posedge		 : VITALDELAYTYPE 	 := 0.72 ns;
	tpw_CLK_negedge		 : VITALDELAYTYPE 	 := 0 ns;
	tperiod_CLK_posedge	 : VITALDELAYTYPE 	 := 1.44 ns;
	tpd_CLK_O		 : VITALDELAYTYPE01Z 	 := (2.74 ns, 2.74 ns, 2.74 ns, 2.74 ns, 2.74 ns, 2.74 ns);
	tpd_OE_O		 : VITALDELAYTYPE01Z 	 := (0.64 ns, 0.64 ns, 0.64 ns, 0.64 ns, 0.64 ns, 0.64 ns)
	);

PORT    (
	O			 : OUT   std_logic;
	D			 : IN    std_logic := 'U';
	CLK			 : IN    std_logic := 'U';
	OE			 : IN    std_logic := 'U'
	);

ATTRIBUTE VITAL_LEVEL0 OF ROT : ENTITY IS TRUE ;

END ROT;
-----------------------------------------------------------------------------
-- ARCHITECTURE declaration
-----------------------------------------------------------------------------
ARCHITECTURE VITAL_VF OF ROT  IS
	ATTRIBUTE VITAL_LEVEL1 OF VITAL_VF : ARCHITECTURE IS TRUE;

	SIGNAL	D_ipd			 : std_ulogic        := 'X';
	SIGNAL	CLK_ipd			 : std_ulogic        := 'X';
	SIGNAL	OE_ipd			 : std_ulogic        := 'X';
	SIGNAL	CLK_dly			 : std_ulogic        := 'X';
	SIGNAL	D_dly			 : std_ulogic        := 'X';
BEGIN
-----------------------------------------------------------------------------
-- INPUT PATH DELAYs
-----------------------------------------------------------------------------
WIREDELAY : BLOCK
BEGIN
	VitalWireDelay( D_ipd, D, tipd_D );
	VitalWireDelay( CLK_ipd, CLK, tipd_CLK );
	VitalWireDelay( OE_ipd, OE, tipd_OE );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
	VitalSignalDelay ( CLK_dly, CLK_ipd, ticd_CLK);
	VitalSignalDelay ( D_dly, D_ipd, tisd_D_CLK);
END BLOCK;

-----------------------------------------------------------------------------
-- Behavior Section
-----------------------------------------------------------------------------
VitalBehaviour_1 : PROCESS(OE_ipd,D_dly,CLK_dly)

VARIABLE 	Tviol_CLK_D_flag1	 : std_ulogic		 := '0';
VARIABLE 	TimingData_D_CLK1	 : VitalTimingDataType	 := VitalTimingDataInit;
VARIABLE 	Tviol_CLK_flag2		 : std_ulogic		 := '0';
VARIABLE 	PeriodData_CLK2		 : VitalPeriodDataType	 := VitalPeriodDataInit;
VARIABLE 	Tviol_CLK_flag3		 : std_ulogic		 := '0';
VARIABLE 	PeriodData_CLK3		 : VitalPeriodDataType	 := VitalPeriodDataInit;
VARIABLE 	Q_int_zd		 : std_ulogic;
VARIABLE 	VCC_zd			 : std_ulogic;
VARIABLE 	PrevDataIn0		 : std_logic_vector (0 to 3) ;
VARIABLE 	O_zd			 : std_ulogic;
VARIABLE 	OGLITCH_DATA		 : VitalGlitchDataType;
VARIABLE 	Violation_Flag		 : std_ulogic;


BEGIN

--Timing Check Section

IF(TimingChecksOn) THEN
VitalSetupHoldCheck(Violation => Tviol_CLK_D_flag1,
TimingData => TimingData_D_CLK1,
TestSignal => D_dly,
TestSignalName => "D",
TestDelay => tisd_D_CLK,
RefSignal => CLK_dly,
RefSignalName => "CLK",
RefDelay => ticd_CLK,
SetupHigh => tsetup_D_CLK_noedge_posedge,
SetupLow => tsetup_D_CLK_noedge_posedge,
HoldHigh => thold_D_CLK_noedge_posedge,
HoldLow => thold_D_CLK_noedge_posedge,
CheckEnabled => ( To_X01( OE_ipd )= '1' ),
RefTransition => '/',
HeaderMsg => InstancePath & "/ROT",
Xon => Xon,
MsgOn => MsgOn,
MsgSeverity => WARNING);

VitalPeriodPulseCheck(Violation => Tviol_CLK_flag2,
PeriodData => PeriodData_CLK2,
TestSignal => CLK_dly,
TestSignalName => "CLK",
TestDelay => ticd_CLK,
Period => 0 ns,
PulseWidthHigh => tpw_CLK_posedge,
PulseWidthLow => tpw_CLK_negedge,
CheckEnabled => ( To_X01( OE_ipd )= '1' ),
HeaderMsg => InstancePath & "/ROT",
Xon => Xon,
MsgOn => MsgOn,
MsgSeverity => WARNING);

VitalPeriodPulseCheck(Violation => Tviol_CLK_flag3,
PeriodData => PeriodData_CLK3,
TestSignal => CLK_dly,
TestSignalName => "CLK",
TestDelay => ticd_CLK,
Period => tperiod_CLK_posedge,
PulseWidthHigh => 0 ns,
PulseWidthLow => 0 ns,
CheckEnabled => posedge( CLK_dly'LAST_VALUE, CLK_dly ) AND ( To_X01( OE_ipd )= '1' ),
HeaderMsg => InstancePath & "/ROT",
Xon => Xon,
MsgOn => MsgOn,
MsgSeverity => WARNING);

END IF;   -- Timing Check Section

--Functionality Section

Violation_Flag	 := ((Tviol_CLK_D_flag1 or Tviol_CLK_flag2) or Tviol_CLK_flag3);
VCC_zd		 := '1';
VitalStateTable(
StateTable => dfftab,
DataIn => std_logic_vector'(D_dly,CLK_dly,VCC_zd,VCC_zd),
Result => Q_int_zd	,
PreviousDataIn => PrevDataIn0);

Q_int_zd	 := (Violation_Flag xor Q_int_zd);
O_zd		 := VitalBUFIF1(Q_int_zd,OE_ipd);

--PathDelay Section

 VitalPathDelay01Z ( O, OGLITCH_DATA, "O", O_zd,
	Paths => (
	0 => ( CLK_dly'LAST_EVENT, tpd_CLK_O, TRUE ),
	1 => ( OE_ipd'LAST_EVENT, tpd_OE_O, TRUE ) ),
	DefaultDelay=>VitalZeroDelay01Z,
	Mode=>VitalInertial,
	XON=>TRUE,
	MsgOn=>TRUE,
	MsgSeverity=>WARNING );


END PROCESS VitalBehaviour_1;
END VITAL_VF;
configuration CFG_ROT_VITAL of ROT is 
        for VITAL_VF
        end for; 
end CFG_ROT_VITAL;
----- VITAL model for cell ROTR -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;

LIBRARY VF1 ;
use VF1.VLOGTOVITAL_TABLES.all;



-- entity declaration --
entity ROTR is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_R_O                        :	VitalDelayType01 := (2.740 ns, 2.740 ns);
      tpd_OE_O                       :	VitalDelayType01z := (0.640 ns, 0.640 ns, 0.640 ns, 0.640 ns, 0.640 ns, 0.640 ns);
      tpd_CLK_O                      :	VitalDelayType01 := (2.740 ns, 2.740 ns);
      tsetup_D_CLK_noedge_posedge :	VitalDelayType := 0.360 ns;
      thold_D_CLK_noedge_posedge :	VitalDelayType := 0.560 ns;
      trecovery_R_CLK_posedge_posedge :	VitalDelayType := 0.330 ns;
      thold_R_CLK_posedge_posedge :	VitalDelayType := 0.530 ns;
      tpw_CLK_posedge :	VitalDelayType := 0.720 ns;
      tperiod_CLK_posedge  :	VitalDelayType := 1.440 ns;
      ticd_CLK                       :	VitalDelayType := 0.000 ns;
      tisd_D_CLK                     :	VitalDelayType := 0.000 ns;
      tisd_R_CLK                     :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_OE                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_R                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      OE                             :	in    STD_ULOGIC;
      R                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      O                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of ROTR : entity is TRUE;
end ROTR;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library VF1;
architecture VITAL_VF of ROTR is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL OE_ipd	 : STD_ULOGIC := 'X';
   SIGNAL R_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL D_CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL R_CLK_dly	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (OE_ipd, OE, tipd_OE);
   VitalWireDelay (R_ipd, R, tipd_R);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   VitalSignalDelay (CLK_dly, CLK_ipd, ticd_CLK);
   VitalSignalDelay (D_CLK_dly, D_ipd, tisd_D_CLK);
   VitalSignalDelay (R_CLK_dly, R_ipd, tisd_R_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (OE_ipd, CLK_dly, D_CLK_dly, R_CLK_dly)

   -- timing check results
   VARIABLE Tviol_D_CLK_OE_EQ_1_AN_R_EQ_1_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_OE_EQ_1_AN_R_EQ_1_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_R_CLK_OE_EQ_1_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_R_CLK_OE_EQ_1_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK_OE_EQ_1_AN_R_EQ_1	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK_OE_EQ_1_AN_R_EQ_1	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_O : STD_LOGIC_VECTOR(0 to 3);
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS O_zdi : STD_LOGIC is Results(1);
   VARIABLE O_zd : STD_ULOGIC := 'X';

   -- output glitch detection variables
   VARIABLE O_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_OE_EQ_1_AN_R_EQ_1_posedge,
          TimingData              => Tmkr_D_CLK_OE_EQ_1_AN_R_EQ_1_posedge,
          TestSignal              => D_CLK_dly,
          TestSignalName          => "D",
          TestDelay               => tisd_D_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          SetupHigh               => tsetup_D_CLK_noedge_posedge,
          SetupLow                => tsetup_D_CLK_noedge_posedge,
          HoldHigh                => thold_D_CLK_noedge_posedge,
          HoldLow                 => thold_D_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT(R_CLK_dly)) AND (OE_ipd)) = '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/ROTR",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_R_CLK_OE_EQ_1_posedge,
          TimingData              => Tmkr_R_CLK_OE_EQ_1_posedge,
          TestSignal              => R_CLK_dly,
          TestSignalName          => "R",
          TestDelay               => tisd_R_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          Recovery                => trecovery_R_CLK_posedge_posedge,
          Removal                 => thold_R_CLK_posedge_posedge,
          ActiveLow               => FALSE,
          CheckEnabled            => 
                           TO_X01(OE_ipd) = '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/ROTR",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK_OE_EQ_1_AN_R_EQ_1,
          PeriodData              => PInfo_CLK_OE_EQ_1_AN_R_EQ_1,
          TestSignal              => CLK_dly,
          TestSignalName          => "CLK",
          TestDelay               => ticd_CLK,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TO_X01((NOT(R_CLK_dly)) AND (OE_ipd)) = '1',
          HeaderMsg               => InstancePath & "/ROTR",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_OE_EQ_1_AN_R_EQ_1_posedge or Tviol_R_CLK_OE_EQ_1_posedge or Pviol_CLK_OE_EQ_1_AN_R_EQ_1;
      VitalStateTable(
        Result => O_zdi,
        PreviousDataIn => PrevData_O,
        StateTable => dfftab,
        DataIn => (
               D_CLK_dly,CLK_dly, NOT(R_CLK_dly),'1'));
      O_zdi := Violation xor O_zdi;
      O_zd := VitalBUFIF1 (O_zdi,OE_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01Z (
       OutSignal => O,
       GlitchData => O_GlitchData,
       OutSignalName => "O",
       OutTemp => O_zd,
       Paths => (0 => (R_CLK_dly'last_event, VitalExtendToFillDelay(tpd_R_O), TRUE),
                 1 => (OE_ipd'last_event, VitalExtendToFillDelay(tpd_OE_O), TRUE),
                 2 => (CLK_dly'last_event, VitalExtendToFillDelay(tpd_CLK_O), TRUE)),
       Mode => VitalInertial,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING,
       OutputMap => "UX01ZWLH-");

end process;
end VITAL_VF;

configuration CFG_ROTR_VITAL of ROTR is 
        for VITAL_VF
        end for; 
end CFG_ROTR_VITAL;
----- VITAL model for cell ROTS -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;

LIBRARY VF1 ;
use VF1.VLOGTOVITAL_TABLES.all;



-- entity declaration --
entity ROTS is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_S_O                        :	VitalDelayType01 := (2.740 ns, 2.740 ns);
      tpd_OE_O                       :	VitalDelayType01z := (0.640 ns, 0.640 ns, 0.640 ns, 0.640 ns, 0.640 ns, 0.640 ns);
      tpd_CLK_O                      :	VitalDelayType01 := (2.740 ns, 2.740 ns);
      tsetup_D_CLK_noedge_posedge :	VitalDelayType := 0.360 ns;
      thold_D_CLK_noedge_posedge :	VitalDelayType := 0.560 ns;
      trecovery_S_CLK_posedge_posedge :	VitalDelayType := 0.330 ns;
      thold_S_CLK_posedge_posedge :	VitalDelayType := 0.530 ns;
      tpw_CLK_posedge :	VitalDelayType := 0.720 ns;
      tperiod_CLK_posedge  :	VitalDelayType := 1.440 ns;
      ticd_CLK                       :	VitalDelayType := 0.000 ns;
      tisd_D_CLK                     :	VitalDelayType := 0.000 ns;
      tisd_S_CLK                     :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_OE                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      OE                             :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      O                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of ROTS : entity is TRUE;
end ROTS;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library VF1;
architecture VITAL_VF of ROTS is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL OE_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL D_CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL S_CLK_dly	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (OE_ipd, OE, tipd_OE);
   VitalWireDelay (S_ipd, S, tipd_S);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   VitalSignalDelay (CLK_dly, CLK_ipd, ticd_CLK);
   VitalSignalDelay (D_CLK_dly, D_ipd, tisd_D_CLK);
   VitalSignalDelay (S_CLK_dly, S_ipd, tisd_S_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (OE_ipd, CLK_dly, D_CLK_dly, S_CLK_dly)

   -- timing check results
   VARIABLE Tviol_D_CLK_OE_EQ_1_AN_S_EQ_1_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_OE_EQ_1_AN_S_EQ_1_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S_CLK_OE_EQ_1_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S_CLK_OE_EQ_1_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK_OE_EQ_1_AN_S_EQ_1	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK_OE_EQ_1_AN_S_EQ_1	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_O : STD_LOGIC_VECTOR(0 to 3);
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS O_zdi : STD_LOGIC is Results(1);
   VARIABLE O_zd : STD_ULOGIC := 'X';

   -- output glitch detection variables
   VARIABLE O_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_OE_EQ_1_AN_S_EQ_1_posedge,
          TimingData              => Tmkr_D_CLK_OE_EQ_1_AN_S_EQ_1_posedge,
          TestSignal              => D_CLK_dly,
          TestSignalName          => "D",
          TestDelay               => tisd_D_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          SetupHigh               => tsetup_D_CLK_noedge_posedge,
          SetupLow                => tsetup_D_CLK_noedge_posedge,
          HoldHigh                => thold_D_CLK_noedge_posedge,
          HoldLow                 => thold_D_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT(S_CLK_dly)) AND (OE_ipd)) = '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/ROTS",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_S_CLK_OE_EQ_1_posedge,
          TimingData              => Tmkr_S_CLK_OE_EQ_1_posedge,
          TestSignal              => S_CLK_dly,
          TestSignalName          => "S",
          TestDelay               => tisd_S_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          Recovery                => trecovery_S_CLK_posedge_posedge,
          Removal                 => thold_S_CLK_posedge_posedge,
          ActiveLow               => FALSE,
          CheckEnabled            => 
                           TO_X01(OE_ipd) = '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/ROTS",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK_OE_EQ_1_AN_S_EQ_1,
          PeriodData              => PInfo_CLK_OE_EQ_1_AN_S_EQ_1,
          TestSignal              => CLK_dly,
          TestSignalName          => "CLK",
          TestDelay               => ticd_CLK,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TO_X01((NOT(S_CLK_dly)) AND (OE_ipd)) = '1',
          HeaderMsg               => InstancePath & "/ROTS",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_OE_EQ_1_AN_S_EQ_1_posedge or Tviol_S_CLK_OE_EQ_1_posedge or Pviol_CLK_OE_EQ_1_AN_S_EQ_1;
      VitalStateTable(
        Result => O_zdi,
        PreviousDataIn => PrevData_O,
        StateTable => dfftab,
        DataIn => (
               D_CLK_dly, CLK_dly, '1',NOT(S_CLK_dly)));
      O_zdi := Violation XOR O_zdi;
      O_zd := VitalBUFIF1 (O_zdi,OE_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01Z (
       OutSignal => O,
       GlitchData => O_GlitchData,
       OutSignalName => "O",
       OutTemp => O_zd,
       Paths => (0 => (S_CLK_dly'last_event, VitalExtendToFillDelay(tpd_S_O), TRUE),
                 1 => (OE_ipd'last_event, VitalExtendToFillDelay(tpd_OE_O), TRUE),
                 2 => (CLK_dly'last_event, VitalExtendToFillDelay(tpd_CLK_O), TRUE)),
       Mode => VitalInertial,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING,
       OutputMap => "UX01ZWLH-");

end process;
end VITAL_VF;

configuration CFG_ROTS_VITAL of ROTS is 
        for VITAL_VF
        end for; 
end CFG_ROTS_VITAL;
----- VITAL model for cell RSFF -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;

LIBRARY VF1 ;
use VF1.VLOGTOVITAL_TABLES.all;



-- entity declaration --
entity RSFF is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_CLK_Q                      :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tsetup_RE_CLK_noedge_posedge   :	VitalDelayType := 2.200 ns;
      thold_RE_CLK_noedge_posedge    :	VitalDelayType := 2.200 ns;
      tsetup_SE_CLK_noedge_posedge   :	VitalDelayType := 2.200 ns;
      thold_SE_CLK_noedge_posedge    :	VitalDelayType := 2.200 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 8.800 ns;
      tpw_CLK_posedge                :	VitalDelayType := 4.400 ns;
      ticd_CLK                       :	VitalDelayType := 0.000 ns;
      tisd_RE_CLK                    :	VitalDelayType := 0.000 ns;
      tisd_SE_CLK                    :	VitalDelayType := 0.000 ns;
      tipd_RE                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_SE                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      RE                             :	in    STD_ULOGIC;
      SE                             :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of RSFF : entity is TRUE;
end RSFF;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library VF1;
architecture VITAL_VF of RSFF is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL RE_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SE_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL RE_CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL SE_CLK_dly	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (RE_ipd, RE, tipd_RE);
   VitalWireDelay (SE_ipd, SE, tipd_SE);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   VitalSignalDelay (CLK_dly, CLK_ipd, ticd_CLK);
   VitalSignalDelay (RE_CLK_dly, RE_ipd, tisd_RE_CLK);
   VitalSignalDelay (SE_CLK_dly, SE_ipd, tisd_SE_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (CLK_dly, RE_CLK_dly, SE_CLK_dly)

   -- timing check results
   VARIABLE Tviol_RE_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_RE_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SE_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SE_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 4);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_RE_CLK_posedge,
          TimingData              => Tmkr_RE_CLK_posedge,
          TestSignal              => RE_CLK_dly,
          TestSignalName          => "RE",
          TestDelay               => tisd_RE_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          SetupHigh               => tsetup_RE_CLK_noedge_posedge,
          SetupLow                => tsetup_RE_CLK_noedge_posedge,
          HoldHigh                => thold_RE_CLK_noedge_posedge,
          HoldLow                 => thold_RE_CLK_noedge_posedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/RSFF",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_SE_CLK_posedge,
          TimingData              => Tmkr_SE_CLK_posedge,
          TestSignal              => SE_CLK_dly,
          TestSignalName          => "SE",
          TestDelay               => tisd_SE_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          SetupHigh               => tsetup_SE_CLK_noedge_posedge,
          SetupLow                => tsetup_SE_CLK_noedge_posedge,
          HoldHigh                => thold_SE_CLK_noedge_posedge,
          HoldLow                 => thold_SE_CLK_noedge_posedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/RSFF",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_dly,
          TestSignalName          => "CLK",
          TestDelay               => ticd_CLK,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/RSFF",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_RE_CLK_posedge or Tviol_SE_CLK_posedge or Pviol_CLK;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => rsfftab,
        DataIn => (
               CLK_dly,RE_CLK_dly,SE_CLK_dly,'1','1'));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (CLK_dly'last_event, tpd_CLK_Q, TRUE)),
       Mode => VitalInertial,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;

configuration CFG_RSFF_VITAL of RSFF is 
        for VITAL_VF
        end for; 
end CFG_RSFF_VITAL;
----- VITAL model for cell RSFFR -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;

LIBRARY VF1 ;
use VF1.VLOGTOVITAL_TABLES.all;



-- entity declaration --
entity RSFFR is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_R_Q                        :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tsetup_RE_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      thold_RE_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      tsetup_SE_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      thold_SE_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      trecovery_R_CLK_posedge_posedge :	VitalDelayType := 2.200 ns;
      thold_R_CLK_posedge_posedge    :	VitalDelayType := 2.200 ns;
      tpw_CLK_posedge         :	VitalDelayType := 4.400 ns;
      tperiod_CLK_posedge             :	VitalDelayType := 8.800 ns;
      ticd_CLK                       :	VitalDelayType := 0.000 ns;
      tisd_RE_CLK                    :	VitalDelayType := 0.000 ns;
      tisd_SE_CLK                    :	VitalDelayType := 0.000 ns;
      tisd_R_CLK                     :	VitalDelayType := 0.000 ns;
      tipd_RE                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_SE                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_R                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      RE                             :	in    STD_ULOGIC;
      SE                             :	in    STD_ULOGIC;
      R                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of RSFFR : entity is TRUE;
end RSFFR;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library VF1;
architecture VITAL_VF of RSFFR is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL RE_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SE_ipd	 : STD_ULOGIC := 'X';
   SIGNAL R_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL RE_CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL SE_CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL R_CLK_dly	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (RE_ipd, RE, tipd_RE);
   VitalWireDelay (SE_ipd, SE, tipd_SE);
   VitalWireDelay (R_ipd, R, tipd_R);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   VitalSignalDelay (CLK_dly, CLK_ipd, ticd_CLK);
   VitalSignalDelay (RE_CLK_dly, RE_ipd, tisd_RE_CLK);
   VitalSignalDelay (SE_CLK_dly, SE_ipd, tisd_SE_CLK);
   VitalSignalDelay (R_CLK_dly, R_ipd, tisd_R_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (CLK_dly, RE_CLK_dly, SE_CLK_dly, R_CLK_dly)

   -- timing check results
   VARIABLE Tviol_RE_CLK_R_EQ_1_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_RE_CLK_R_EQ_1_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SE_CLK_R_EQ_1_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SE_CLK_R_EQ_1_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_R_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_R_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK_R_EQ_1	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK_R_EQ_1	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 4);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_RE_CLK_R_EQ_1_posedge,
          TimingData              => Tmkr_RE_CLK_R_EQ_1_posedge,
          TestSignal              => RE_CLK_dly,
          TestSignalName          => "RE",
          TestDelay               => tisd_RE_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          SetupHigh               => tsetup_RE_CLK_noedge_posedge,
          SetupLow                => tsetup_RE_CLK_noedge_posedge,
          HoldHigh                => thold_RE_CLK_noedge_posedge,
          HoldLow                 => thold_RE_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(R_CLK_dly) = '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/RSFFR",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_SE_CLK_R_EQ_1_posedge,
          TimingData              => Tmkr_SE_CLK_R_EQ_1_posedge,
          TestSignal              => SE_CLK_dly,
          TestSignalName          => "SE",
          TestDelay               => tisd_SE_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          SetupHigh               => tsetup_SE_CLK_noedge_posedge,
          SetupLow                => tsetup_SE_CLK_noedge_posedge,
          HoldHigh                => thold_SE_CLK_noedge_posedge,
          HoldLow                 => thold_SE_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(R_CLK_dly) = '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/RSFFR",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_R_CLK_posedge,
          TimingData              => Tmkr_R_CLK_posedge,
          TestSignal              => R_CLK_dly,
          TestSignalName          => "R",
          TestDelay               => tisd_R_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          Recovery                => trecovery_R_CLK_posedge_posedge,
          Removal                 => thold_R_CLK_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/RSFFR",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK_R_EQ_1,
          PeriodData              => PInfo_CLK_R_EQ_1,
          TestSignal              => CLK_dly,
          TestSignalName          => "CLK",
          TestDelay               => ticd_CLK,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TO_X01((R_CLK_dly) ) = '1',
          HeaderMsg               => InstancePath & "/RSFFR",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_RE_CLK_R_EQ_1_posedge or Tviol_SE_CLK_R_EQ_1_posedge or Pviol_CLK_R_EQ_1 or Tviol_R_CLK_posedge;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => rsfftab,
        DataIn => (
                CLK_dly, RE_CLK_dly, SE_CLK_dly, '1', R_CLK_dly));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (R_CLK_dly'last_event, tpd_R_Q, TRUE),
                 1 => (CLK_dly'last_event, tpd_CLK_Q, TRUE)),
       Mode => VitalInertial,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;

configuration CFG_RSFFR_VITAL of RSFFR is 
        for VITAL_VF
        end for; 
end CFG_RSFFR_VITAL;
----- VITAL model for cell RSFFRH -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;

LIBRARY VF1 ;
use VF1.VLOGTOVITAL_TABLES.all;



-- entity declaration --
entity RSFFRH is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_R_Q                        :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tsetup_RE_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      thold_RE_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      tsetup_SE_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      thold_SE_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      trecovery_R_CLK_negedge_posedge :	VitalDelayType := 2.200 ns;
      thold_R_CLK_negedge_posedge    :	VitalDelayType := 2.200 ns;
      tpw_CLK_posedge         :	VitalDelayType := 4.400 ns;
      tpw_R_posedge         :	VitalDelayType := 4.400 ns;
      tperiod_CLK_posedge             :	VitalDelayType := 8.800 ns;
      ticd_CLK                       :	VitalDelayType := 0.000 ns;
      tisd_RE_CLK                    :	VitalDelayType := 0.000 ns;
      tisd_SE_CLK                    :	VitalDelayType := 0.000 ns;
      tisd_R_CLK                     :	VitalDelayType := 0.000 ns;
      tipd_RE                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_SE                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_R                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      RE                             :	in    STD_ULOGIC;
      SE                             :	in    STD_ULOGIC;
      R                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of RSFFRH : entity is TRUE;
end RSFFRH;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library VF1;
architecture VITAL_VF of RSFFRH is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL RE_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SE_ipd	 : STD_ULOGIC := 'X';
   SIGNAL R_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL RE_CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL SE_CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL R_CLK_dly	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (RE_ipd, RE, tipd_RE);
   VitalWireDelay (SE_ipd, SE, tipd_SE);
   VitalWireDelay (R_ipd, R, tipd_R);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   VitalSignalDelay (CLK_dly, CLK_ipd, ticd_CLK);
   VitalSignalDelay (RE_CLK_dly, RE_ipd, tisd_RE_CLK);
   VitalSignalDelay (SE_CLK_dly, SE_ipd, tisd_SE_CLK);
   VitalSignalDelay (R_CLK_dly, R_ipd, tisd_R_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (CLK_dly, RE_CLK_dly, SE_CLK_dly, R_CLK_dly)

   -- timing check results
   VARIABLE Tviol_RE_CLK_R_EQ_0_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_RE_CLK_R_EQ_0_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SE_CLK_R_EQ_0_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SE_CLK_R_EQ_0_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_R_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_R_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK_R_EQ_0	: STD_ULOGIC := '0';
   VARIABLE Pviol_R	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK_R_EQ_0	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE PInfo_R	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 4);
   VARIABLE R_inverted : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_RE_CLK_R_EQ_0_posedge,
          TimingData              => Tmkr_RE_CLK_R_EQ_0_posedge,
          TestSignal              => RE_CLK_dly,
          TestSignalName          => "RE",
          TestDelay               => tisd_RE_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          SetupHigh               => tsetup_RE_CLK_noedge_posedge,
          SetupLow                => tsetup_RE_CLK_noedge_posedge,
          HoldHigh                => thold_RE_CLK_noedge_posedge,
          HoldLow                 => thold_RE_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(R_CLK_dly) = '0',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/RSFFRH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_SE_CLK_R_EQ_0_posedge,
          TimingData              => Tmkr_SE_CLK_R_EQ_0_posedge,
          TestSignal              => SE_CLK_dly,
          TestSignalName          => "SE",
          TestDelay               => tisd_SE_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          SetupHigh               => tsetup_SE_CLK_noedge_posedge,
          SetupLow                => tsetup_SE_CLK_noedge_posedge,
          HoldHigh                => thold_SE_CLK_noedge_posedge,
          HoldLow                 => thold_SE_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(R_CLK_dly) = '0',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/RSFFRH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_R_CLK_posedge,
          TimingData              => Tmkr_R_CLK_posedge,
          TestSignal              => R_CLK_dly,
          TestSignalName          => "R",
          TestDelay               => tisd_R_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          Recovery                => trecovery_R_CLK_negedge_posedge,
          Removal                 => thold_R_CLK_negedge_posedge,
          ActiveLow               => FALSE,
          CheckEnabled            => TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/RSFFRH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_R,
          PeriodData              => PInfo_R,
          TestSignal              => R_CLK_dly,
          TestSignalName          => "R",
          TestDelay               => tisd_R_CLK,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_R_posedge,
          CheckEnabled            => TRUE, 
          HeaderMsg               => InstancePath & "/RSFFRH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK_R_EQ_0,
          PeriodData              => PInfo_CLK_R_EQ_0,
          TestSignal              => CLK_dly,
          TestSignalName          => "CLK",
          TestDelay               => ticd_CLK,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TO_X01(R_CLK_dly ) = '0',
          HeaderMsg               => InstancePath & "/RSFFRH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_RE_CLK_R_EQ_0_posedge or Tviol_R_CLK_posedge or Pviol_CLK_R_EQ_0 or Tviol_SE_CLK_R_EQ_0_posedge or Pviol_R;
      R_inverted := (NOT R_CLK_dly);
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => rsfftab,
        DataIn => (
               CLK_dly, RE_CLK_dly, SE_CLK_dly, '1', R_inverted));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (R_CLK_dly'last_event, tpd_R_Q, TRUE),
                 1 => (CLK_dly'last_event, tpd_CLK_Q, TRUE)),
       Mode => VitalInertial,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;

configuration CFG_RSFFRH_VITAL of RSFFRH is 
        for VITAL_VF
        end for; 
end CFG_RSFFRH_VITAL;
----- VITAL model for cell RSFFRS -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;
library VF1;
use VF1.VLOGTOVITAL_TABLES.all;


-- entity declaration --
entity RSFFRS is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_R_Q                        :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tpd_S_Q                        :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tsetup_RE_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      thold_RE_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      tsetup_SE_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      thold_SE_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      trecovery_R_CLK_posedge_posedge :	VitalDelayType := 2.200 ns;
      thold_R_CLK_posedge_posedge :	VitalDelayType := 2.200 ns;
      trecovery_S_CLK_posedge_posedge :	VitalDelayType := 2.200 ns;
      thold_S_CLK_posedge_posedge :	VitalDelayType := 2.200 ns;
      tpw_CLK_posedge :	VitalDelayType := 4.400 ns;
      tpw_R_negedge :	VitalDelayType := 4.400 ns;
      tpw_S_negedge :	VitalDelayType := 4.400 ns;
      tperiod_CLK_posedge   :	VitalDelayType := 8.800 ns;
      ticd_CLK                       :	VitalDelayType := 0.000 ns;
      tisd_RE_CLK                    :	VitalDelayType := 0.000 ns;
      tisd_SE_CLK                    :	VitalDelayType := 0.000 ns;
      tisd_R_CLK                     :	VitalDelayType := 0.000 ns;
      tisd_S_CLK                     :	VitalDelayType := 0.000 ns;
      tipd_RE                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_SE                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_R                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      RE                             :	in    STD_ULOGIC;
      SE                             :	in    STD_ULOGIC;
      R                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of RSFFRS : entity is TRUE;
end RSFFRS;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library VF1;
use VF1.VLOGTOVITAL_TABLES.all;
architecture VITAL_VF of RSFFRS is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL RE_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SE_ipd	 : STD_ULOGIC := 'X';
   SIGNAL R_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL RE_CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL SE_CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL R_CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL S_CLK_dly	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (RE_ipd, RE, tipd_RE);
   VitalWireDelay (SE_ipd, SE, tipd_SE);
   VitalWireDelay (R_ipd, R, tipd_R);
   VitalWireDelay (S_ipd, S, tipd_S);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   VitalSignalDelay (CLK_dly, CLK_ipd, ticd_CLK);
   VitalSignalDelay (RE_CLK_dly, RE_ipd, tisd_RE_CLK);
   VitalSignalDelay (SE_CLK_dly, SE_ipd, tisd_SE_CLK);
   VitalSignalDelay (R_CLK_dly, R_ipd, tisd_R_CLK);
   VitalSignalDelay (S_CLK_dly, S_ipd, tisd_S_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (CLK_dly, RE_CLK_dly, SE_CLK_dly, R_CLK_dly, S_CLK_dly)

   -- timing check results
   VARIABLE Tviol_RE_CLK_R_EQ_1_AN_S_EQ_1_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_RE_CLK_R_EQ_1_AN_S_EQ_1_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SE_CLK_R_EQ_1_AN_S_EQ_1_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SE_CLK_R_EQ_1_AN_S_EQ_1_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_R_CLK_S_EQ_1_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_R_CLK_S_EQ_1_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S_CLK_R_EQ_1_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S_CLK_R_EQ_1_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK_R_EQ_1_AN_S_EQ_1	: STD_ULOGIC := '0';
   VARIABLE Pviol_R	: STD_ULOGIC := '0';
   VARIABLE Pviol_S	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK_R_EQ_1_AN_S_EQ_1	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE PInfo_R	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE PInfo_S	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(1 to 5);
   VARIABLE RE_delayed : STD_ULOGIC := 'X';
   VARIABLE SE_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_RE_CLK_R_EQ_1_AN_S_EQ_1_posedge,
          TimingData              => Tmkr_RE_CLK_R_EQ_1_AN_S_EQ_1_posedge,
          TestSignal              => RE_CLK_dly,
          TestSignalName          => "RE",
          TestDelay               => tisd_RE_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          SetupHigh               => tsetup_RE_CLK_noedge_posedge,
          SetupLow                => tsetup_RE_CLK_noedge_posedge,
          HoldHigh                => thold_RE_CLK_noedge_posedge,
          HoldLow                 => thold_RE_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((S_CLK_dly) AND (R_CLK_dly)) /= '0',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/RSFFRS",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_SE_CLK_R_EQ_1_AN_S_EQ_1_posedge,
          TimingData              => Tmkr_SE_CLK_R_EQ_1_AN_S_EQ_1_posedge,
          TestSignal              => SE_CLK_dly,
          TestSignalName          => "SE",
          TestDelay               => tisd_SE_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          SetupHigh               => tsetup_SE_CLK_noedge_posedge,
          SetupLow                => tsetup_SE_CLK_noedge_posedge,
          HoldHigh                => thold_SE_CLK_noedge_posedge,
          HoldLow                 => thold_SE_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((S_CLK_dly) AND (R_CLK_dly)) /= '0',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/RSFFRS",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_R_CLK_S_EQ_1_posedge,
          TimingData              => Tmkr_R_CLK_S_EQ_1_posedge,
          TestSignal              => R_CLK_dly,
          TestSignalName          => "R",
          TestDelay               => tisd_R_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          Recovery                => trecovery_R_CLK_posedge_posedge,
          Removal                 => thold_R_CLK_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TO_X01(S_CLK_dly) /= '0',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/RSFFRS",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_S_CLK_R_EQ_1_posedge,
          TimingData              => Tmkr_S_CLK_R_EQ_1_posedge,
          TestSignal              => S_CLK_dly,
          TestSignalName          => "S",
          TestDelay               => tisd_S_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          Recovery                => trecovery_S_CLK_posedge_posedge,
          Removal                 => thold_S_CLK_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TO_X01(R_CLK_dly) /= '0',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/RSFFRS",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_S,
          PeriodData              => PInfo_S,
          TestSignal              => S_CLK_dly,
          TestSignalName          => "S",
          TestDelay               => tisd_S_CLK,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_S_negedge,
          CheckEnabled            => TRUE, 
          HeaderMsg               => InstancePath & "/RSFFRS",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_R,
          PeriodData              => PInfo_R,
          TestSignal              => R_CLK_dly,
          TestSignalName          => "R",
          TestDelay               => tisd_R_CLK,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_R_negedge,
          CheckEnabled            => TRUE, 
          HeaderMsg               => InstancePath & "/RSFFRS",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK_R_EQ_1_AN_S_EQ_1,
          PeriodData              => PInfo_CLK_R_EQ_1_AN_S_EQ_1,
          TestSignal              => CLK_dly,
          TestSignalName          => "CLK",
          TestDelay               => ticd_CLK,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TO_X01(( (NOT S_CLK_dly) ) OR ( (NOT R_CLK_dly) )
                            ) /= '1',
          HeaderMsg               => InstancePath & "/RSFFRS",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_RE_CLK_R_EQ_1_AN_S_EQ_1_posedge or Tviol_R_CLK_S_EQ_1_posedge or Tviol_SE_CLK_R_EQ_1_AN_S_EQ_1_posedge or Tviol_S_CLK_R_EQ_1_posedge or Pviol_CLK_R_EQ_1_AN_S_EQ_1 or Pviol_R or Pviol_S ;
      --VitalStateTable(
       -- Result => QBAR_zd,
        --PreviousDataIn => PrevData_QBAR,
        --StateTable => RSFFRS_QBAR_tab,
        --DataIn => (
         --      S_CLK_dly, CLK_delayed, RE_delayed, SE_delayed, Q_zd, R_CLK_dly, CLK_dly));
      --QBAR_zd := Violation XOR QBAR_zd;
      RE_delayed := RE_CLK_dly;
      SE_delayed := SE_CLK_dly;
      CLK_delayed := CLK_dly;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => rsfftab,
        DataIn => (
               CLK_dly, RE_delayed, SE_delayed, S_CLK_dly, R_CLK_dly));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (R_CLK_dly'last_event, tpd_R_Q, TRUE),
                 1 => (S_CLK_dly'last_event, tpd_S_Q, TRUE),
                 2 => (CLK_dly'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;

configuration CFG_RSFFRS_VITAL of RSFFRS is 
        for VITAL_VF
        end for; 
end CFG_RSFFRS_VITAL;
----- VITAL model for cell RSFFRSH -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;
library VF1;
use VF1.VLOGTOVITAL_TABLES.all;


-- entity declaration --
entity RSFFRSH is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_R_Q                        :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tpd_S_Q                        :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tsetup_RE_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      thold_RE_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      tsetup_SE_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      thold_SE_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      trecovery_R_CLK_negedge_posedge :	VitalDelayType := 2.200 ns;
      thold_R_CLK_negedge_posedge :	VitalDelayType := 2.200 ns;
      trecovery_S_CLK_negedge_posedge :	VitalDelayType := 2.200 ns;
      thold_S_CLK_negedge_posedge :	VitalDelayType := 2.200 ns;
      tpw_CLK_posedge :	VitalDelayType := 4.400 ns;
      tpw_R_posedge :	VitalDelayType := 4.400 ns;
      tpw_S_posedge :	VitalDelayType := 4.400 ns;
      tperiod_CLK_posedge   :	VitalDelayType := 8.800 ns;
      ticd_CLK                       :	VitalDelayType := 0.000 ns;
      tisd_RE_CLK                    :	VitalDelayType := 0.000 ns;
      tisd_SE_CLK                    :	VitalDelayType := 0.000 ns;
      tisd_R_CLK                     :	VitalDelayType := 0.000 ns;
      tisd_S_CLK                     :	VitalDelayType := 0.000 ns;
      tipd_RE                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_SE                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_R                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      RE                             :	in    STD_ULOGIC;
      SE                             :	in    STD_ULOGIC;
      R                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of RSFFRSH : entity is TRUE;
end RSFFRSH;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library VF1;
use VF1.VLOGTOVITAL_TABLES.all;
architecture VITAL_VF of RSFFRSH is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL RE_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SE_ipd	 : STD_ULOGIC := 'X';
   SIGNAL R_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL RE_CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL SE_CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL R_CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL S_CLK_dly	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (RE_ipd, RE, tipd_RE);
   VitalWireDelay (SE_ipd, SE, tipd_SE);
   VitalWireDelay (R_ipd, R, tipd_R);
   VitalWireDelay (S_ipd, S, tipd_S);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   VitalSignalDelay (CLK_dly, CLK_ipd, ticd_CLK);
   VitalSignalDelay (RE_CLK_dly, RE_ipd, tisd_RE_CLK);
   VitalSignalDelay (SE_CLK_dly, SE_ipd, tisd_SE_CLK);
   VitalSignalDelay (R_CLK_dly, R_ipd, tisd_R_CLK);
   VitalSignalDelay (S_CLK_dly, S_ipd, tisd_S_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (CLK_dly, RE_CLK_dly, SE_CLK_dly, R_CLK_dly, S_CLK_dly)

   -- timing check results
   VARIABLE Tviol_RE_CLK_R_EQ_0_AN_S_EQ_0_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_RE_CLK_R_EQ_0_AN_S_EQ_0_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SE_CLK_R_EQ_0_AN_S_EQ_0_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SE_CLK_R_EQ_0_AN_S_EQ_0_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_R_CLK_S_EQ_0_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_R_CLK_S_EQ_0_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S_CLK_R_EQ_0_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S_CLK_R_EQ_0_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK_R_EQ_0_AN_S_EQ_0	: STD_ULOGIC := '0';
   VARIABLE Pviol_R	: STD_ULOGIC := '0';
   VARIABLE Pviol_S	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK_R_EQ_0_AN_S_EQ_0	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE PInfo_R	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE PInfo_S	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(1 to 5);
   VARIABLE R_inverted : STD_ULOGIC := 'X';
   VARIABLE S_inverted : STD_ULOGIC := 'X';
   VARIABLE RE_delayed : STD_ULOGIC := 'X';
   VARIABLE SE_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_RE_CLK_R_EQ_0_AN_S_EQ_0_posedge,
          TimingData              => Tmkr_RE_CLK_R_EQ_0_AN_S_EQ_0_posedge,
          TestSignal              => RE_CLK_dly,
          TestSignalName          => "RE",
          TestDelay               => tisd_RE_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          SetupHigh               => tsetup_RE_CLK_noedge_posedge,
          SetupLow                => tsetup_RE_CLK_noedge_posedge,
          HoldHigh                => thold_RE_CLK_noedge_posedge,
          HoldLow                 => thold_RE_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(((NOT S_CLK_dly)) AND ((NOT R_CLK_dly))) /=
                            '0',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/RSFFRSH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_SE_CLK_R_EQ_0_AN_S_EQ_0_posedge,
          TimingData              => Tmkr_SE_CLK_R_EQ_0_AN_S_EQ_0_posedge,
          TestSignal              => SE_CLK_dly,
          TestSignalName          => "SE",
          TestDelay               => tisd_SE_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          SetupHigh               => tsetup_SE_CLK_noedge_posedge,
          SetupLow                => tsetup_SE_CLK_noedge_posedge,
          HoldHigh                => thold_SE_CLK_noedge_posedge,
          HoldLow                 => thold_SE_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(((NOT S_CLK_dly)) AND ((NOT R_CLK_dly))) /=
                            '0',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/RSFFRSH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_R_CLK_S_EQ_0_posedge,
          TimingData              => Tmkr_R_CLK_S_EQ_0_posedge,
          TestSignal              => R_CLK_dly,
          TestSignalName          => "R",
          TestDelay               => tisd_R_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          Recovery                => trecovery_R_CLK_negedge_posedge,
          Removal                 => thold_R_CLK_negedge_posedge,
          ActiveLow               => FALSE,
          CheckEnabled            => 
                           TO_X01((NOT S_CLK_dly)) /= '0',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/RSFFRSH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_S_CLK_R_EQ_0_posedge,
          TimingData              => Tmkr_S_CLK_R_EQ_0_posedge,
          TestSignal              => S_CLK_dly,
          TestSignalName          => "S",
          TestDelay               => tisd_S_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          Recovery                => trecovery_S_CLK_negedge_posedge,
          Removal                 => thold_S_CLK_negedge_posedge,
          ActiveLow               => FALSE,
          CheckEnabled            => 
                           TO_X01((NOT R_CLK_dly)) /= '0',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/RSFFRSH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_S,
          PeriodData              => PInfo_S,
          TestSignal              => S_CLK_dly,
          TestSignalName          => "S",
          TestDelay               => tisd_S_CLK,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_S_posedge,
          CheckEnabled            => TRUE, 
          HeaderMsg               => InstancePath & "/RSFFRSH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_R,
          PeriodData              => PInfo_R,
          TestSignal              => R_CLK_dly,
          TestSignalName          => "R",
          TestDelay               => tisd_R_CLK,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_R_posedge,
          CheckEnabled            => TRUE, 
          HeaderMsg               => InstancePath & "/RSFFRSH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK_R_EQ_0_AN_S_EQ_0,
          PeriodData              => PInfo_CLK_R_EQ_0_AN_S_EQ_0,
          TestSignal              => CLK_dly,
          TestSignalName          => "CLK",
          TestDelay               => ticd_CLK,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TO_X01(( S_CLK_dly ) OR ( R_CLK_dly ) ) /= '1',
          HeaderMsg               => InstancePath & "/RSFFRSH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_RE_CLK_R_EQ_0_AN_S_EQ_0_posedge or Tviol_SE_CLK_R_EQ_0_AN_S_EQ_0_posedge or Tviol_S_CLK_R_EQ_0_posedge or Pviol_CLK_R_EQ_0_AN_S_EQ_0 or Tviol_R_CLK_S_EQ_0_posedge or Pviol_R or Pviol_S;
      R_inverted := NOT R_CLK_dly;
      S_inverted := NOT S_CLK_dly;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => rsfftab,
        DataIn => (
               CLK_dly, RE_CLK_dly, SE_CLK_dly, S_inverted, R_inverted));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (R_CLK_dly'last_event, tpd_R_Q, TRUE),
                 1 => (S_CLK_dly'last_event, tpd_S_Q, TRUE),
                 2 => (CLK_dly'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;

configuration CFG_RSFFRSH_VITAL of RSFFRSH is 
        for VITAL_VF
        end for; 
end CFG_RSFFRSH_VITAL;
----- VITAL model for cell RSFFRSS -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;

LIBRARY VF1 ;
use VF1.VLOGTOVITAL_TABLES.all;



-- entity declaration --
entity RSFFRSS is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_R_Q                        :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tpd_S_Q                        :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tsetup_RE_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      thold_RE_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      tsetup_SE_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      thold_SE_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      trecovery_R_CLK_negedge_posedge :	VitalDelayType := 2.200 ns;
      thold_R_CLK_negedge_posedge :	VitalDelayType := 2.200 ns;
      trecovery_S_CLK_negedge_posedge :	VitalDelayType := 2.200 ns;
      thold_S_CLK_negedge_posedge :	VitalDelayType := 2.200 ns;
      tpw_CLK_posedge :	VitalDelayType := 4.400 ns;
      tperiod_CLK_posedge  :	VitalDelayType := 8.800 ns;
      ticd_CLK                       :	VitalDelayType := 0.000 ns;
      tisd_RE_CLK                    :	VitalDelayType := 0.000 ns;
      tisd_SE_CLK                    :	VitalDelayType := 0.000 ns;
      tisd_R_CLK                     :	VitalDelayType := 0.000 ns;
      tisd_S_CLK                     :	VitalDelayType := 0.000 ns;
      tipd_RE                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_SE                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_R                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      RE                             :	in    STD_ULOGIC;
      SE                             :	in    STD_ULOGIC;
      R                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of RSFFRSS : entity is TRUE;
end RSFFRSS;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library VF1;
architecture VITAL_VF of RSFFRSS is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL RE_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SE_ipd	 : STD_ULOGIC := 'X';
   SIGNAL R_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL RE_CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL SE_CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL R_CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL S_CLK_dly	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (RE_ipd, RE, tipd_RE);
   VitalWireDelay (SE_ipd, SE, tipd_SE);
   VitalWireDelay (R_ipd, R, tipd_R);
   VitalWireDelay (S_ipd, S, tipd_S);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   VitalSignalDelay (CLK_dly, CLK_ipd, ticd_CLK);
   VitalSignalDelay (RE_CLK_dly, RE_ipd, tisd_RE_CLK);
   VitalSignalDelay (SE_CLK_dly, SE_ipd, tisd_SE_CLK);
   VitalSignalDelay (R_CLK_dly, R_ipd, tisd_R_CLK);
   VitalSignalDelay (S_CLK_dly, S_ipd, tisd_S_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (CLK_dly, RE_CLK_dly, SE_CLK_dly, R_CLK_dly, S_CLK_dly)

   -- timing check results
   VARIABLE Tviol_RE_CLK_R_EQ_0_ANB_S_EQ_0_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_RE_CLK_R_EQ_0_ANB_S_EQ_0_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SE_CLK_R_EQ_0_ANB_S_EQ_0_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SE_CLK_R_EQ_0_ANB_S_EQ_0_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_R_CLK_S_EQ_0_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_R_CLK_S_EQ_0_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S_CLK_R_EQ_0_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S_CLK_R_EQ_0_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK_R_EQ_0_ANB_S_EQ_0	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK_R_EQ_0_ANB_S_EQ_0	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 4);
   VARIABLE R_inverted : STD_ULOGIC := 'X';
   VARIABLE S_inverted : STD_ULOGIC := 'X';
   VARIABLE RE_in : STD_ULOGIC := 'X';
   VARIABLE SE_in : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_RE_CLK_R_EQ_0_ANB_S_EQ_0_posedge,
          TimingData              => Tmkr_RE_CLK_R_EQ_0_ANB_S_EQ_0_posedge,
          TestSignal              => RE_CLK_dly,
          TestSignalName          => "RE",
          TestDelay               => tisd_RE_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          SetupHigh               => tsetup_RE_CLK_noedge_posedge,
          SetupLow                => tsetup_RE_CLK_noedge_posedge,
          HoldHigh                => thold_RE_CLK_noedge_posedge,
          HoldLow                 => thold_RE_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(((NOT S_CLK_dly)) AND ((NOT R_CLK_dly))) = '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/RSFFRSS",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_SE_CLK_R_EQ_0_ANB_S_EQ_0_posedge,
          TimingData              => Tmkr_SE_CLK_R_EQ_0_ANB_S_EQ_0_posedge,
          TestSignal              => SE_CLK_dly,
          TestSignalName          => "SE",
          TestDelay               => tisd_SE_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          SetupHigh               => tsetup_SE_CLK_noedge_posedge,
          SetupLow                => tsetup_SE_CLK_noedge_posedge,
          HoldHigh                => thold_SE_CLK_noedge_posedge,
          HoldLow                 => thold_SE_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(((NOT S_CLK_dly)) AND ((NOT R_CLK_dly))) = '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/RSFFRSS",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_R_CLK_S_EQ_0_posedge,
          TimingData              => Tmkr_R_CLK_S_EQ_0_posedge,
          TestSignal              => R_CLK_dly,
          TestSignalName          => "R",
          TestDelay               => tisd_R_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          Recovery                => trecovery_R_CLK_negedge_posedge,
          Removal                 => thold_R_CLK_negedge_posedge,
          ActiveLow               => FALSE,
          CheckEnabled            => 
                           TO_X01((S_CLK_dly)) = '0',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/RSFFRSS",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_S_CLK_R_EQ_0_posedge,
          TimingData              => Tmkr_S_CLK_R_EQ_0_posedge,
          TestSignal              => S_CLK_dly,
          TestSignalName          => "S",
          TestDelay               => tisd_S_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          Recovery                => trecovery_S_CLK_negedge_posedge,
          Removal                 => thold_S_CLK_negedge_posedge,
          ActiveLow               => FALSE,
          CheckEnabled            => 
                           TO_X01((R_CLK_dly)) = '0',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/RSFFRSS",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK_R_EQ_0_ANB_S_EQ_0,
          PeriodData              => PInfo_CLK_R_EQ_0_ANB_S_EQ_0,
          TestSignal              => CLK_dly,
          TestSignalName          => "CLK",
          TestDelay               => ticd_CLK,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TO_X01(( NOT S_CLK_dly ) AND ( NOT R_CLK_dly ) ) = '1',
          HeaderMsg               => InstancePath & "/RSFFRSS",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_RE_CLK_R_EQ_0_ANB_S_EQ_0_posedge or Tviol_SE_CLK_R_EQ_0_ANB_S_EQ_0_posedge or Tviol_R_CLK_S_EQ_0_posedge or Tviol_S_CLK_R_EQ_0_posedge or Pviol_CLK_R_EQ_0_ANB_S_EQ_0;
      R_inverted := (NOT R_CLK_dly);
      S_inverted := (NOT S_CLK_dly);
      SE_in := VitalOR2 (S_inverted,SE_CLK_dly);
      RE_in := VitalAND2 (S_CLK_dly,RE_CLK_dly);
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => rsfftab,
        DataIn => (
               CLK_dly, RE_in, SE_in, '1', R_CLK_dly));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (R_CLK_dly'last_event, tpd_R_Q, TRUE),
                 1 => (S_CLK_dly'last_event, tpd_S_Q, TRUE),
                 2 => (CLK_dly'last_event, tpd_CLK_Q, TRUE)),
       Mode => VitalInertial,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;

configuration CFG_RSFFRSS_VITAL of RSFFRSS is 
        for VITAL_VF
        end for; 
end CFG_RSFFRSS_VITAL;

----------------------------------------------------------------
-- 
-- Created by the Synopsys Library Compiler v3.4a
-- FILENAME     :    VF1_VITAL.vhd
-- FILE CONTENTS:    Entity, Structural Architecture(VITAL),
--                   and Configuration
-- DATE CREATED :    Tue Jun 10 12:17:07 1997
-- 
-- LIBRARY      :    VF1
-- REVISION     :    Not Specified
-- TECHNOLOGY   :    cmos
-- TIME SCALE   :    1 ns
-- LOGIC SYSTEM :    IEEE-1164
-- NOTES        :    VITAL, TimingChecksOn(TRUE), XGenerationOn(TRUE), TimingMessage(TRUE), VitalInertial 
-- HISTORY      :
-- 
----------------------------------------------------------------

----- VITAL model for cell RSFFRSSH -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;

LIBRARY VF1 ;
use VF1.VLOGTOVITAL_TABLES.all;



-- entity declaration --
entity RSFFRSSH is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_R_Q                        :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tpd_S_Q                        :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tsetup_RE_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      thold_RE_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      tsetup_SE_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      thold_SE_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      trecovery_R_CLK_negedge_posedge :	VitalDelayType := 2.200 ns;
      thold_R_CLK_negedge_posedge :	VitalDelayType := 2.200 ns;
      tsetup_S_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      thold_S_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      tpw_CLK_posedge :	VitalDelayType := 4.400 ns;
      tpw_R_posedge :	VitalDelayType := 4.400 ns;
      tperiod_CLK_posedge  :	VitalDelayType := 8.800 ns;
      ticd_CLK                       :	VitalDelayType := 0.000 ns;
      tisd_RE_CLK                    :	VitalDelayType := 0.000 ns;
      tisd_SE_CLK                    :	VitalDelayType := 0.000 ns;
      tisd_R_CLK                     :	VitalDelayType := 0.000 ns;
      tisd_S_CLK                     :	VitalDelayType := 0.000 ns;
      tipd_RE                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_SE                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_R                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      RE                             :	in    STD_ULOGIC;
      SE                             :	in    STD_ULOGIC;
      R                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of RSFFRSSH : entity is TRUE;
end RSFFRSSH;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library VF1;
architecture VITAL_VF of RSFFRSSH is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL RE_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SE_ipd	 : STD_ULOGIC := 'X';
   SIGNAL R_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL RE_CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL SE_CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL R_CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL S_CLK_dly	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (RE_ipd, RE, tipd_RE);
   VitalWireDelay (SE_ipd, SE, tipd_SE);
   VitalWireDelay (R_ipd, R, tipd_R);
   VitalWireDelay (S_ipd, S, tipd_S);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   VitalSignalDelay (CLK_dly, CLK_ipd, ticd_CLK);
   VitalSignalDelay (RE_CLK_dly, RE_ipd, tisd_RE_CLK);
   VitalSignalDelay (SE_CLK_dly, SE_ipd, tisd_SE_CLK);
   VitalSignalDelay (R_CLK_dly, R_ipd, tisd_R_CLK);
   VitalSignalDelay (S_CLK_dly, S_ipd, tisd_S_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (CLK_dly, RE_CLK_dly, SE_CLK_dly, R_CLK_dly, S_CLK_dly)

   -- timing check results
   VARIABLE Tviol_RE_CLK_R_EQ_0_ANB_S_EQ_0_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_RE_CLK_R_EQ_0_ANB_S_EQ_0_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SE_CLK_R_EQ_0_ANB_S_EQ_0_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SE_CLK_R_EQ_0_ANB_S_EQ_0_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_R_CLK_S_EQ_0_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_R_CLK_S_EQ_0_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S_CLK_R_EQ_0_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S_CLK_R_EQ_0_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK_R_EQ_0_ANB_S_EQ_0	: STD_ULOGIC := '0';
   VARIABLE Pviol_R	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK_R_EQ_0_ANB_S_EQ_0	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE PInfo_R	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 4);
   VARIABLE R_inverted : STD_ULOGIC := 'X';
   VARIABLE S_inverted : STD_ULOGIC := 'X';
   VARIABLE RE_in : STD_ULOGIC := 'X';
   VARIABLE SE_in : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_RE_CLK_R_EQ_0_ANB_S_EQ_0_posedge,
          TimingData              => Tmkr_RE_CLK_R_EQ_0_ANB_S_EQ_0_posedge,
          TestSignal              => RE_CLK_dly,
          TestSignalName          => "RE",
          TestDelay               => tisd_RE_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          SetupHigh               => tsetup_RE_CLK_noedge_posedge,
          SetupLow                => tsetup_RE_CLK_noedge_posedge,
          HoldHigh                => thold_RE_CLK_noedge_posedge,
          HoldLow                 => thold_RE_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(((NOT S_CLK_dly)) AND ((NOT R_CLK_dly))) = '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/RSFFRSSH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_SE_CLK_R_EQ_0_ANB_S_EQ_0_posedge,
          TimingData              => Tmkr_SE_CLK_R_EQ_0_ANB_S_EQ_0_posedge,
          TestSignal              => SE_CLK_dly,
          TestSignalName          => "SE",
          TestDelay               => tisd_SE_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          SetupHigh               => tsetup_SE_CLK_noedge_posedge,
          SetupLow                => tsetup_SE_CLK_noedge_posedge,
          HoldHigh                => thold_SE_CLK_noedge_posedge,
          HoldLow                 => thold_SE_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(((NOT S_CLK_dly)) AND ((NOT R_CLK_dly))) = '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/RSFFRSSH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_R_CLK_S_EQ_0_posedge,
          TimingData              => Tmkr_R_CLK_S_EQ_0_posedge,
          TestSignal              => R_CLK_dly,
          TestSignalName          => "R",
          TestDelay               => tisd_R_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          Recovery                => trecovery_R_CLK_negedge_posedge,
          Removal                 => thold_R_CLK_negedge_posedge,
          ActiveLow               => FALSE,
          CheckEnabled            => 
                           TO_X01((S_CLK_dly)) = '0',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/RSFFRSSH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_S_CLK_R_EQ_0_posedge,
          TimingData              => Tmkr_S_CLK_R_EQ_0_posedge,
          TestSignal              => S_CLK_dly,
          TestSignalName          => "S",
          TestDelay               => tisd_S_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          SetupHigh               => tsetup_S_CLK_noedge_posedge,
          SetupLow                => tsetup_S_CLK_noedge_posedge,
          HoldHigh                => thold_S_CLK_noedge_posedge,
          HoldLow                 => thold_S_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((R_CLK_dly)) = '0',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/RSFFRSSH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_R,
          PeriodData              => PInfo_R,
          TestSignal              => R_CLK_dly,
          TestSignalName          => "R",
          TestDelay               => tisd_R_CLK,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_R_posedge,
          CheckEnabled            => TRUE, 
          HeaderMsg               => InstancePath & "/RSFFRSSH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK_R_EQ_0_ANB_S_EQ_0,
          PeriodData              => PInfo_CLK_R_EQ_0_ANB_S_EQ_0,
          TestSignal              => CLK_dly,
          TestSignalName          => "CLK",
          TestDelay               => ticd_CLK,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TO_X01(( NOT S_CLK_dly ) AND ( NOT R_CLK_dly ) ) = '1',
          HeaderMsg               => InstancePath & "/RSFFRSSH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_RE_CLK_R_EQ_0_ANB_S_EQ_0_posedge or Tviol_SE_CLK_R_EQ_0_ANB_S_EQ_0_posedge or Tviol_R_CLK_S_EQ_0_posedge or Tviol_S_CLK_R_EQ_0_posedge or Pviol_CLK_R_EQ_0_ANB_S_EQ_0 or Pviol_R;
      R_inverted := (NOT R_CLK_dly);
      S_inverted := (NOT S_CLK_dly);
      RE_in := VitalAND2 (S_inverted,RE_CLK_dly);
      SE_in := VitalOR2 (S_CLK_dly,SE_CLK_dly);
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => rsfftab,
        DataIn => (
               CLK_dly, RE_in, SE_in, '1', R_inverted));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (R_CLK_dly'last_event, tpd_R_Q, TRUE),
                 1 => (S_CLK_dly'last_event, tpd_S_Q, TRUE),
                 2 => (CLK_dly'last_event, tpd_CLK_Q, TRUE)),
       Mode => VitalInertial,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_VF;
configuration CFG_RSFFRSSH_VITAL of RSFFRSSH is 
        for VITAL_VF
        end for; 
end CFG_RSFFRSSH_VITAL;
----- VITAL model for cell RSFFS -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;

LIBRARY VF1 ;
use VF1.VLOGTOVITAL_TABLES.all;



-- entity declaration --
entity RSFFS is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_S_Q                        :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tsetup_RE_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      thold_RE_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      tsetup_SE_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      thold_SE_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      trecovery_S_CLK_posedge_posedge :	VitalDelayType := 2.200 ns;
      thold_S_CLK_posedge_posedge    :	VitalDelayType := 2.200 ns;
      tpw_CLK_posedge         :	VitalDelayType := 4.400 ns;
      tperiod_CLK_posedge             :	VitalDelayType := 8.800 ns;
      ticd_CLK                       :	VitalDelayType := 0.000 ns;
      tisd_RE_CLK                    :	VitalDelayType := 0.000 ns;
      tisd_SE_CLK                    :	VitalDelayType := 0.000 ns;
      tisd_S_CLK                     :	VitalDelayType := 0.000 ns;
      tipd_RE                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_SE                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      RE                             :	in    STD_ULOGIC;
      SE                             :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of RSFFS : entity is TRUE;
end RSFFS;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library VF1;
architecture VITAL_VF of RSFFS is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL RE_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SE_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL RE_CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL SE_CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL S_CLK_dly	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (RE_ipd, RE, tipd_RE);
   VitalWireDelay (SE_ipd, SE, tipd_SE);
   VitalWireDelay (S_ipd, S, tipd_S);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   VitalSignalDelay (CLK_dly, CLK_ipd, ticd_CLK);
   VitalSignalDelay (RE_CLK_dly, RE_ipd, tisd_RE_CLK);
   VitalSignalDelay (SE_CLK_dly, SE_ipd, tisd_SE_CLK);
   VitalSignalDelay (S_CLK_dly, S_ipd, tisd_S_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (CLK_dly, RE_CLK_dly, SE_CLK_dly, S_CLK_dly)

   -- timing check results
   VARIABLE Tviol_RE_CLK_S_EQ_1_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_RE_CLK_S_EQ_1_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SE_CLK_S_EQ_1_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SE_CLK_S_EQ_1_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK_S_EQ_1	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK_S_EQ_1	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 4);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_RE_CLK_S_EQ_1_posedge,
          TimingData              => Tmkr_RE_CLK_S_EQ_1_posedge,
          TestSignal              => RE_CLK_dly,
          TestSignalName          => "RE",
          TestDelay               => tisd_RE_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          SetupHigh               => tsetup_RE_CLK_noedge_posedge,
          SetupLow                => tsetup_RE_CLK_noedge_posedge,
          HoldHigh                => thold_RE_CLK_noedge_posedge,
          HoldLow                 => thold_RE_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(S_CLK_dly) = '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/RSFFS",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_SE_CLK_S_EQ_1_posedge,
          TimingData              => Tmkr_SE_CLK_S_EQ_1_posedge,
          TestSignal              => SE_CLK_dly,
          TestSignalName          => "SE",
          TestDelay               => tisd_SE_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          SetupHigh               => tsetup_SE_CLK_noedge_posedge,
          SetupLow                => tsetup_SE_CLK_noedge_posedge,
          HoldHigh                => thold_SE_CLK_noedge_posedge,
          HoldLow                 => thold_SE_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(S_CLK_dly) = '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/RSFFS",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_S_CLK_posedge,
          TimingData              => Tmkr_S_CLK_posedge,
          TestSignal              => S_CLK_dly,
          TestSignalName          => "S",
          TestDelay               => tisd_S_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          Recovery                => trecovery_S_CLK_posedge_posedge,
          Removal                 => thold_S_CLK_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/RSFFS",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK_S_EQ_1,
          PeriodData              => PInfo_CLK_S_EQ_1,
          TestSignal              => CLK_dly,
          TestSignalName          => "CLK",
          TestDelay               => ticd_CLK,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TO_X01((S_CLK_dly) ) = '1',
          HeaderMsg               => InstancePath & "/RSFFS",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_RE_CLK_S_EQ_1_posedge or Tviol_S_CLK_posedge or Pviol_CLK_S_EQ_1 or Tviol_SE_CLK_S_EQ_1_posedge;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => rsfftab,
        DataIn => (
               CLK_dly, RE_CLK_dly, SE_CLK_dly, S_CLK_dly, '1'));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (S_CLK_dly'last_event, tpd_S_Q, TRUE),
                 1 => (CLK_dly'last_event, tpd_CLK_Q, TRUE)),
       Mode => VitalInertial,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;

configuration CFG_RSFFS_VITAL of RSFFS is 
        for VITAL_VF
        end for; 
end CFG_RSFFS_VITAL;
----- VITAL model for cell RSFFSH -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;

LIBRARY VF1 ;
use VF1.VLOGTOVITAL_TABLES.all;



-- entity declaration --
entity RSFFSH is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_S_Q                        :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tsetup_RE_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      thold_RE_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      tsetup_SE_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      thold_SE_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      trecovery_S_CLK_negedge_posedge :	VitalDelayType := 2.200 ns;
      thold_S_CLK_negedge_posedge    :	VitalDelayType := 2.200 ns;
      tpw_CLK_posedge         :	VitalDelayType := 4.400 ns;
      tpw_S_posedge         :	VitalDelayType := 4.400 ns;
      tperiod_CLK_posedge             :	VitalDelayType := 8.800 ns;
      ticd_CLK                       :	VitalDelayType := 0.000 ns;
      tisd_RE_CLK                    :	VitalDelayType := 0.000 ns;
      tisd_SE_CLK                    :	VitalDelayType := 0.000 ns;
      tisd_S_CLK                     :	VitalDelayType := 0.000 ns;
      tipd_RE                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_SE                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      RE                             :	in    STD_ULOGIC;
      SE                             :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of RSFFSH : entity is TRUE;
end RSFFSH;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library VF1;
architecture VITAL_VF of RSFFSH is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL RE_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SE_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL RE_CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL SE_CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL S_CLK_dly	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (RE_ipd, RE, tipd_RE);
   VitalWireDelay (SE_ipd, SE, tipd_SE);
   VitalWireDelay (S_ipd, S, tipd_S);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   VitalSignalDelay (CLK_dly, CLK_ipd, ticd_CLK);
   VitalSignalDelay (RE_CLK_dly, RE_ipd, tisd_RE_CLK);
   VitalSignalDelay (SE_CLK_dly, SE_ipd, tisd_SE_CLK);
   VitalSignalDelay (S_CLK_dly, S_ipd, tisd_S_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (CLK_dly, RE_CLK_dly, SE_CLK_dly, S_CLK_dly)

   -- timing check results
   VARIABLE Tviol_RE_CLK_S_EQ_0_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_RE_CLK_S_EQ_0_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SE_CLK_S_EQ_0_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SE_CLK_S_EQ_0_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK_S_EQ_0	: STD_ULOGIC := '0';
   VARIABLE Pviol_S	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK_S_EQ_0	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE PInfo_S	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 4);
   VARIABLE S_inverted : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_RE_CLK_S_EQ_0_posedge,
          TimingData              => Tmkr_RE_CLK_S_EQ_0_posedge,
          TestSignal              => RE_CLK_dly,
          TestSignalName          => "RE",
          TestDelay               => tisd_RE_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          SetupHigh               => tsetup_RE_CLK_noedge_posedge,
          SetupLow                => tsetup_RE_CLK_noedge_posedge,
          HoldHigh                => thold_RE_CLK_noedge_posedge,
          HoldLow                 => thold_RE_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(S_CLK_dly) = '0',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/RSFFSH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_SE_CLK_S_EQ_0_posedge,
          TimingData              => Tmkr_SE_CLK_S_EQ_0_posedge,
          TestSignal              => SE_CLK_dly,
          TestSignalName          => "SE",
          TestDelay               => tisd_SE_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          SetupHigh               => tsetup_SE_CLK_noedge_posedge,
          SetupLow                => tsetup_SE_CLK_noedge_posedge,
          HoldHigh                => thold_SE_CLK_noedge_posedge,
          HoldLow                 => thold_SE_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(S_CLK_dly) = '0',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/RSFFSH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_S_CLK_posedge,
          TimingData              => Tmkr_S_CLK_posedge,
          TestSignal              => S_CLK_dly,
          TestSignalName          => "S",
          TestDelay               => tisd_S_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          Recovery                => trecovery_S_CLK_negedge_posedge,
          Removal                 => thold_S_CLK_negedge_posedge,
          ActiveLow               => FALSE,
          CheckEnabled            => TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/RSFFSH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_S,
          PeriodData              => PInfo_S,
          TestSignal              => S_CLK_dly,
          TestSignalName          => "S",
          TestDelay               => tisd_S_CLK,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_S_posedge,
          CheckEnabled            => TRUE, 
          HeaderMsg               => InstancePath & "/RSFFSH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK_S_EQ_0,
          PeriodData              => PInfo_CLK_S_EQ_0,
          TestSignal              => CLK_dly,
          TestSignalName          => "CLK",
          TestDelay               => ticd_CLK,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TO_X01(S_CLK_dly ) = '0',
          HeaderMsg               => InstancePath & "/RSFFSH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_RE_CLK_S_EQ_0_posedge or Tviol_S_CLK_posedge or Tviol_SE_CLK_S_EQ_0_posedge or Pviol_CLK_S_EQ_0;
      S_inverted := (NOT S_CLK_dly);
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => rsfftab,
        DataIn => (
               CLK_dly, RE_CLK_dly, SE_CLK_dly, S_inverted, '1'));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (S_CLK_dly'last_event, tpd_S_Q, TRUE),
                 1 => (CLK_dly'last_event, tpd_CLK_Q, TRUE)),
       Mode => VitalInertial,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;

configuration CFG_RSFFSH_VITAL of RSFFSH is 
        for VITAL_VF
        end for; 
end CFG_RSFFSH_VITAL;
----- VITAL model for cell TFF -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;

LIBRARY VF1 ;
use VF1.VLOGTOVITAL_TABLES.all;



-- entity declaration --
entity TFF is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_CLK_Q                      :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tsetup_T_CLK_noedge_posedge    :	VitalDelayType := 2.200 ns;
      thold_T_CLK_noedge_posedge     :	VitalDelayType := 2.200 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 8.800 ns;
      tpw_CLK_posedge                :	VitalDelayType := 4.400 ns;
      ticd_CLK                       :	VitalDelayType := 0.000 ns;
      tisd_T_CLK                     :	VitalDelayType := 0.000 ns;
      tipd_T                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      T                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of TFF : entity is TRUE;
end TFF;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library VF1;
architecture VITAL_VF of TFF is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL T_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL T_CLK_dly	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (T_ipd, T, tipd_T);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   VitalSignalDelay (CLK_dly, CLK_ipd, ticd_CLK);
   VitalSignalDelay (T_CLK_dly, T_ipd, tisd_T_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (CLK_dly, T_CLK_dly)

   -- timing check results
   VARIABLE Tviol_T_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_T_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 3);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => '0');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_T_CLK_posedge,
          TimingData              => Tmkr_T_CLK_posedge,
          TestSignal              => T_CLK_dly,
          TestSignalName          => "T",
          TestDelay               => tisd_T_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          SetupHigh               => tsetup_T_CLK_noedge_posedge,
          SetupLow                => tsetup_T_CLK_noedge_posedge,
          HoldHigh                => thold_T_CLK_noedge_posedge,
          HoldLow                 => thold_T_CLK_noedge_posedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/TFF",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_dly,
          TestSignalName          => "CLK",
          TestDelay               => ticd_CLK,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/TFF",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_T_CLK_posedge or Pviol_CLK;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => tfftab,
        DataIn => (
               CLK_dly, T_CLK_dly, '1', '1'));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (CLK_dly'last_event, tpd_CLK_Q, TRUE)),
       Mode => VitalInertial,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;

configuration CFG_TFF_VITAL of TFF is 
        for VITAL_VF
        end for; 
end CFG_TFF_VITAL;
----- VITAL model for cell TFFR -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;

LIBRARY VF1 ;
use VF1.VLOGTOVITAL_TABLES.all;



-- entity declaration --
entity TFFR is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_R_Q                        :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tsetup_T_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      thold_T_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      trecovery_R_CLK_posedge_posedge :	VitalDelayType := 2.200 ns;
      thold_R_CLK_posedge_posedge    :	VitalDelayType := 2.200 ns;
      tpw_CLK_posedge         :	VitalDelayType := 4.400 ns;
      tperiod_CLK_posedge             :	VitalDelayType := 8.800 ns;
      ticd_CLK                       :	VitalDelayType := 0.000 ns;
      tisd_T_CLK                     :	VitalDelayType := 0.000 ns;
      tisd_R_CLK                     :	VitalDelayType := 0.000 ns;
      tipd_T                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_R                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      T                              :	in    STD_ULOGIC;
      R                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of TFFR : entity is TRUE;
end TFFR;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library VF1;
architecture VITAL_VF of TFFR is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL T_ipd	 : STD_ULOGIC := 'X';
   SIGNAL R_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL T_CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL R_CLK_dly	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (T_ipd, T, tipd_T);
   VitalWireDelay (R_ipd, R, tipd_R);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   VitalSignalDelay (CLK_dly, CLK_ipd, ticd_CLK);
   VitalSignalDelay (T_CLK_dly, T_ipd, tisd_T_CLK);
   VitalSignalDelay (R_CLK_dly, R_ipd, tisd_R_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (CLK_dly, T_CLK_dly, R_CLK_dly)

   -- timing check results
   VARIABLE Tviol_T_CLK_R_EQ_1_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_T_CLK_R_EQ_1_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_R_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_R_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK_R_EQ_1	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK_R_EQ_1	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 3);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_T_CLK_R_EQ_1_posedge,
          TimingData              => Tmkr_T_CLK_R_EQ_1_posedge,
          TestSignal              => T_CLK_dly,
          TestSignalName          => "T",
          TestDelay               => tisd_T_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          SetupHigh               => tsetup_T_CLK_noedge_posedge,
          SetupLow                => tsetup_T_CLK_noedge_posedge,
          HoldHigh                => thold_T_CLK_noedge_posedge,
          HoldLow                 => thold_T_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(R_CLK_dly) = '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/TFFR",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_R_CLK_posedge,
          TimingData              => Tmkr_R_CLK_posedge,
          TestSignal              => R_CLK_dly,
          TestSignalName          => "R",
          TestDelay               => tisd_R_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          Recovery                => trecovery_R_CLK_posedge_posedge,
          Removal                 => thold_R_CLK_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/TFFR",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK_R_EQ_1,
          PeriodData              => PInfo_CLK_R_EQ_1,
          TestSignal              => CLK_dly,
          TestSignalName          => "CLK",
          TestDelay               => ticd_CLK,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TO_X01((R_CLK_dly) ) = '1',
          HeaderMsg               => InstancePath & "/TFFR",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_T_CLK_R_EQ_1_posedge or Pviol_CLK_R_EQ_1 or Tviol_R_CLK_posedge;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => tfftab,
        DataIn => (
               CLK_dly, T_CLK_dly, '1', R_CLK_dly));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (R_CLK_dly'last_event, tpd_R_Q, TRUE),
                 1 => (CLK_dly'last_event, tpd_CLK_Q, TRUE)),
       Mode => VitalInertial,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;

configuration CFG_TFFR_VITAL of TFFR is 
        for VITAL_VF
        end for; 
end CFG_TFFR_VITAL;
----- VITAL model for cell TFFRH -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;

LIBRARY VF1 ;
use VF1.VLOGTOVITAL_TABLES.all;



-- entity declaration --
entity TFFRH is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_R_Q                        :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tsetup_T_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      thold_T_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      trecovery_R_CLK_negedge_posedge :	VitalDelayType := 2.200 ns;
      thold_R_CLK_negedge_posedge    :	VitalDelayType := 2.200 ns;
      tpw_CLK_posedge         :	VitalDelayType := 4.400 ns;
      tpw_R_posedge         :	VitalDelayType := 4.400 ns;
      tperiod_CLK_posedge             :	VitalDelayType := 8.800 ns;
      ticd_CLK                       :	VitalDelayType := 0.000 ns;
      tisd_T_CLK                     :	VitalDelayType := 0.000 ns;
      tisd_R_CLK                     :	VitalDelayType := 0.000 ns;
      tipd_T                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_R                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      T                              :	in    STD_ULOGIC;
      R                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of TFFRH : entity is TRUE;
end TFFRH;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library VF1;
architecture VITAL_VF of TFFRH is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL T_ipd	 : STD_ULOGIC := 'X';
   SIGNAL R_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL T_CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL R_CLK_dly	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (T_ipd, T, tipd_T);
   VitalWireDelay (R_ipd, R, tipd_R);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   VitalSignalDelay (CLK_dly, CLK_ipd, ticd_CLK);
   VitalSignalDelay (T_CLK_dly, T_ipd, tisd_T_CLK);
   VitalSignalDelay (R_CLK_dly, R_ipd, tisd_R_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (CLK_dly, T_CLK_dly, R_CLK_dly)

   -- timing check results
   VARIABLE Tviol_T_CLK_R_EQ_0_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_T_CLK_R_EQ_0_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_R_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_R_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK_R_EQ_0	: STD_ULOGIC := '0';
   VARIABLE Pviol_R	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK_R_EQ_0	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE PInfo_R	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 3);
   VARIABLE R_inverted : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_T_CLK_R_EQ_0_posedge,
          TimingData              => Tmkr_T_CLK_R_EQ_0_posedge,
          TestSignal              => T_CLK_dly,
          TestSignalName          => "T",
          TestDelay               => tisd_T_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          SetupHigh               => tsetup_T_CLK_noedge_posedge,
          SetupLow                => tsetup_T_CLK_noedge_posedge,
          HoldHigh                => thold_T_CLK_noedge_posedge,
          HoldLow                 => thold_T_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((R_CLK_dly)) = '0',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/TFFRH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_R_CLK_posedge,
          TimingData              => Tmkr_R_CLK_posedge,
          TestSignal              => R_CLK_dly,
          TestSignalName          => "R",
          TestDelay               => tisd_R_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          Recovery                => trecovery_R_CLK_negedge_posedge,
          Removal                 => thold_R_CLK_negedge_posedge,
          ActiveLow               => FALSE,
          CheckEnabled            => TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/TFFRH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_R,
          PeriodData              => PInfo_R,
          TestSignal              => R_CLK_dly,
          TestSignalName          => "R",
          TestDelay               => tisd_R_CLK,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_R_posedge,
          CheckEnabled            => TRUE, 
          HeaderMsg               => InstancePath & "/TFFRH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK_R_EQ_0,
          PeriodData              => PInfo_CLK_R_EQ_0,
          TestSignal              => CLK_dly,
          TestSignalName          => "CLK",
          TestDelay               => ticd_CLK,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TO_X01(R_CLK_dly ) = '0',
          HeaderMsg               => InstancePath & "/TFFRH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_T_CLK_R_EQ_0_posedge or Tviol_R_CLK_posedge or Pviol_CLK_R_EQ_0;
      R_inverted := (NOT R_CLK_dly);
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => tfftab,
        DataIn => (
               CLK_dly, T_CLK_dly, '1', R_inverted));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (R_CLK_dly'last_event, tpd_R_Q, TRUE),
                 1 => (CLK_dly'last_event, tpd_CLK_Q, TRUE)),
       Mode => VitalInertial,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;

configuration CFG_TFFRH_VITAL of TFFRH is 
        for VITAL_VF
        end for; 
end CFG_TFFRH_VITAL;
----- VITAL model for cell TFFRS -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;
LIBRARY VF1 ;
use VF1.VLOGTOVITAL_TABLES.all;


-- entity declaration --
entity TFFRS is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_S_Q                        :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tpd_R_Q                        :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tsetup_T_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      thold_T_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      trecovery_R_CLK_posedge_posedge :	VitalDelayType := 2.200 ns;
      thold_R_CLK_posedge_posedge :	VitalDelayType := 2.200 ns;
      trecovery_S_CLK_posedge_posedge :	VitalDelayType := 2.200 ns;
      thold_S_CLK_posedge_posedge :	VitalDelayType := 2.200 ns;
      tpw_CLK_posedge :	VitalDelayType := 4.400 ns;
      tpw_R_negedge :	VitalDelayType := 4.400 ns;
      tpw_S_negedge :	VitalDelayType := 4.400 ns;
      tperiod_CLK_posedge   :	VitalDelayType := 8.800 ns;
      ticd_CLK                       :	VitalDelayType := 0.000 ns;
      tisd_T_CLK                     :	VitalDelayType := 0.000 ns;
      tisd_R_CLK                     :	VitalDelayType := 0.000 ns;
      tisd_S_CLK                     :	VitalDelayType := 0.000 ns;
      tipd_T                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_R                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      T                              :	in    STD_ULOGIC;
      R                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of TFFRS : entity is TRUE;
end TFFRS;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library VF1;
architecture VITAL_VF of TFFRS is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL T_ipd	 : STD_ULOGIC := 'X';
   SIGNAL R_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL T_CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL R_CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL S_CLK_dly	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (T_ipd, T, tipd_T);
   VitalWireDelay (R_ipd, R, tipd_R);
   VitalWireDelay (S_ipd, S, tipd_S);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   VitalSignalDelay (CLK_dly, CLK_ipd, ticd_CLK);
   VitalSignalDelay (T_CLK_dly, T_ipd, tisd_T_CLK);
   VitalSignalDelay (R_CLK_dly, R_ipd, tisd_R_CLK);
   VitalSignalDelay (S_CLK_dly, S_ipd, tisd_S_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (CLK_dly, T_CLK_dly, R_CLK_dly, S_CLK_dly)

   -- timing check results
   VARIABLE Tviol_T_CLK_R_EQ_1_AN_S_EQ_1_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_T_CLK_R_EQ_1_AN_S_EQ_1_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_R_CLK_S_EQ_1_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_R_CLK_S_EQ_1_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S_CLK_R_EQ_1_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S_CLK_R_EQ_1_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK_R_EQ_1_AN_S_EQ_1	: STD_ULOGIC := '0';
   VARIABLE Pviol_R	: STD_ULOGIC := '0';
   VARIABLE Pviol_S	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK_R_EQ_1_AN_S_EQ_1	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE PInfo_R	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE PInfo_S	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(1 to 4);
   VARIABLE T_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_T_CLK_R_EQ_1_AN_S_EQ_1_posedge,
          TimingData              => Tmkr_T_CLK_R_EQ_1_AN_S_EQ_1_posedge,
          TestSignal              => T_CLK_dly,
          TestSignalName          => "T",
          TestDelay               => tisd_T_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          SetupHigh               => tsetup_T_CLK_noedge_posedge,
          SetupLow                => tsetup_T_CLK_noedge_posedge,
          HoldHigh                => thold_T_CLK_noedge_posedge,
          HoldLow                 => thold_T_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((S_CLK_dly) AND (R_CLK_dly)) /= '0',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/TFFRS",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_R_CLK_S_EQ_1_posedge,
          TimingData              => Tmkr_R_CLK_S_EQ_1_posedge,
          TestSignal              => R_CLK_dly,
          TestSignalName          => "R",
          TestDelay               => tisd_R_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          Recovery                => trecovery_R_CLK_posedge_posedge,
          Removal                 => thold_R_CLK_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TO_X01(S_CLK_dly) /= '0',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/TFFRS",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_S_CLK_R_EQ_1_posedge,
          TimingData              => Tmkr_S_CLK_R_EQ_1_posedge,
          TestSignal              => S_CLK_dly,
          TestSignalName          => "S",
          TestDelay               => tisd_S_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          Recovery                => trecovery_S_CLK_posedge_posedge,
          Removal                 => thold_S_CLK_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TO_X01(R_CLK_dly) /= '0',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/TFFRS",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_S,
          PeriodData              => PInfo_S,
          TestSignal              => S_CLK_dly,
          TestSignalName          => "S",
          TestDelay               => tisd_S_CLK,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_S_negedge,
          CheckEnabled            => TRUE, 
          HeaderMsg               => InstancePath & "/TFFRS",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_R,
          PeriodData              => PInfo_R,
          TestSignal              => R_CLK_dly,
          TestSignalName          => "R",
          TestDelay               => tisd_R_CLK,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_R_negedge,
          CheckEnabled            => TRUE, 
          HeaderMsg               => InstancePath & "/TFFRS",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK_R_EQ_1_AN_S_EQ_1,
          PeriodData              => PInfo_CLK_R_EQ_1_AN_S_EQ_1,
          TestSignal              => CLK_dly,
          TestSignalName          => "CLK",
          TestDelay               => ticd_CLK,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TO_X01(( (NOT S_CLK_dly) ) OR ( (NOT R_CLK_dly) )
                            ) /= '1',
          HeaderMsg               => InstancePath & "/TFFRS",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_T_CLK_R_EQ_1_AN_S_EQ_1_posedge or Tviol_R_CLK_S_EQ_1_posedge or Tviol_S_CLK_R_EQ_1_posedge or Pviol_CLK_R_EQ_1_AN_S_EQ_1 or Pviol_R or Pviol_s;
      T_delayed := T_CLK_dly;
      CLK_delayed := CLK_dly;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => tfftab,
        DataIn => (
               CLK_dly, T_CLK_dly,S_CLK_dly, R_CLK_dly));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (S_CLK_dly'last_event, tpd_S_Q, TRUE),
                 1 => (R_CLK_dly'last_event, tpd_R_Q, TRUE),
                 2 => (CLK_dly'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;

configuration CFG_TFFRS_VITAL of TFFRS is 
        for VITAL_VF
        end for; 
end CFG_TFFRS_VITAL;
----- VITAL model for cell TFFRSH -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;
LIBRARY VF1 ;
use VF1.VLOGTOVITAL_TABLES.all;

-- entity declaration --
entity TFFRSH is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_S_Q                        :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tpd_R_Q                        :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tsetup_T_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      thold_T_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      trecovery_R_CLK_negedge_posedge :	VitalDelayType := 2.200 ns;
      thold_R_CLK_negedge_posedge :	VitalDelayType := 2.200 ns;
      trecovery_S_CLK_negedge_posedge :	VitalDelayType := 2.200 ns;
      thold_S_CLK_negedge_posedge :	VitalDelayType := 2.200 ns;
      tpw_CLK_posedge :	VitalDelayType := 4.400 ns;
      tpw_R_posedge :	VitalDelayType := 4.400 ns;
      tpw_S_posedge :	VitalDelayType := 4.400 ns;
      tperiod_CLK_posedge   :	VitalDelayType := 8.800 ns;
      ticd_CLK                       :	VitalDelayType := 0.000 ns;
      tisd_T_CLK                     :	VitalDelayType := 0.000 ns;
      tisd_R_CLK                     :	VitalDelayType := 0.000 ns;
      tisd_S_CLK                     :	VitalDelayType := 0.000 ns;
      tipd_T                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_R                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      T                              :	in    STD_ULOGIC;
      R                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of TFFRSH : entity is TRUE;
end TFFRSH;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library VF1;
architecture VITAL_VF of TFFRSH is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL T_ipd	 : STD_ULOGIC := 'X';
   SIGNAL R_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL T_CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL R_CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL S_CLK_dly	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (T_ipd, T, tipd_T);
   VitalWireDelay (R_ipd, R, tipd_R);
   VitalWireDelay (S_ipd, S, tipd_S);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   VitalSignalDelay (CLK_dly, CLK_ipd, ticd_CLK);
   VitalSignalDelay (T_CLK_dly, T_ipd, tisd_T_CLK);
   VitalSignalDelay (R_CLK_dly, R_ipd, tisd_R_CLK);
   VitalSignalDelay (S_CLK_dly, S_ipd, tisd_S_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (CLK_dly, T_CLK_dly, R_CLK_dly, S_CLK_dly)

   -- timing check results
   VARIABLE Tviol_T_CLK_R_EQ_0_AN_S_EQ_0_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_T_CLK_R_EQ_0_AN_S_EQ_0_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_R_CLK_S_EQ_0_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_R_CLK_S_EQ_0_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S_CLK_R_EQ_0_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S_CLK_R_EQ_0_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK_R_EQ_0_AN_S_EQ_0	: STD_ULOGIC := '0';
   VARIABLE Pviol_R	: STD_ULOGIC := '0';
   VARIABLE Pviol_S	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK_R_EQ_0_AN_S_EQ_0	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE PInfo_R	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE PInfo_S	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(1 to 4);
   VARIABLE T_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE S_inverted : STD_ULOGIC := 'X';
   VARIABLE R_inverted : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_T_CLK_R_EQ_0_AN_S_EQ_0_posedge,
          TimingData              => Tmkr_T_CLK_R_EQ_0_AN_S_EQ_0_posedge,
          TestSignal              => T_CLK_dly,
          TestSignalName          => "T",
          TestDelay               => tisd_T_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          SetupHigh               => tsetup_T_CLK_noedge_posedge,
          SetupLow                => tsetup_T_CLK_noedge_posedge,
          HoldHigh                => thold_T_CLK_noedge_posedge,
          HoldLow                 => thold_T_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(((NOT S_CLK_dly)) AND ((NOT R_CLK_dly))) /=
                            '0',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/TFFRSH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_R_CLK_S_EQ_0_posedge,
          TimingData              => Tmkr_R_CLK_S_EQ_0_posedge,
          TestSignal              => R_CLK_dly,
          TestSignalName          => "R",
          TestDelay               => tisd_R_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          Recovery                => trecovery_R_CLK_negedge_posedge,
          Removal                 => thold_R_CLK_negedge_posedge,
          ActiveLow               => FALSE,
          CheckEnabled            => 
                           TO_X01((NOT S_CLK_dly)) /= '0',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/TFFRSH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_S_CLK_R_EQ_0_posedge,
          TimingData              => Tmkr_S_CLK_R_EQ_0_posedge,
          TestSignal              => S_CLK_dly,
          TestSignalName          => "S",
          TestDelay               => tisd_S_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          Recovery                => trecovery_S_CLK_negedge_posedge,
          Removal                 => thold_S_CLK_negedge_posedge,
          ActiveLow               => FALSE,
          CheckEnabled            => 
                           TO_X01((NOT R_CLK_dly)) /= '0',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/TFFRSH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_S,
          PeriodData              => PInfo_S,
          TestSignal              => S_CLK_dly,
          TestSignalName          => "S",
          TestDelay               => tisd_S_CLK,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_S_posedge,
          CheckEnabled            => TRUE, 
          HeaderMsg               => InstancePath & "/TFFRSH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_R,
          PeriodData              => PInfo_R,
          TestSignal              => R_CLK_dly,
          TestSignalName          => "R",
          TestDelay               => tisd_R_CLK,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_R_posedge,
          CheckEnabled            => TRUE, 
          HeaderMsg               => InstancePath & "/TFFRSH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK_R_EQ_0_AN_S_EQ_0,
          PeriodData              => PInfo_CLK_R_EQ_0_AN_S_EQ_0,
          TestSignal              => CLK_dly,
          TestSignalName          => "CLK",
          TestDelay               => ticd_CLK,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TO_X01(( S_CLK_dly ) OR ( R_CLK_dly ) ) /= '1',
          HeaderMsg               => InstancePath & "/TFFRSH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_T_CLK_R_EQ_0_AN_S_EQ_0_posedge or Tviol_S_CLK_R_EQ_0_posedge or Pviol_CLK_R_EQ_0_AN_S_EQ_0 or Tviol_R_CLK_S_EQ_0_posedge or Pviol_R or Pviol_S;
      T_delayed := T_CLK_dly;
      CLK_delayed := CLK_dly;
      S_inverted := NOT S_CLK_dly;
      R_inverted := NOT R_CLK_dly;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => tfftab,
        DataIn => (
               CLK_dly, T_CLK_dly,S_inverted, R_inverted));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (S_CLK_dly'last_event, tpd_S_Q, TRUE),
                 1 => (R_CLK_dly'last_event, tpd_R_Q, TRUE),
                 2 => (CLK_dly'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;

configuration CFG_TFFRSH_VITAL of TFFRSH is 
        for VITAL_VF
        end for; 
end CFG_TFFRSH_VITAL;
----- VITAL model for cell TFFRSS -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;

LIBRARY VF1 ;
use VF1.VLOGTOVITAL_TABLES.all;



-- entity declaration --
entity TFFRSS is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_S_Q                        :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tpd_R_Q                        :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tsetup_T_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      thold_T_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      trecovery_R_CLK_posedge_posedge :	VitalDelayType := 2.200 ns;
      thold_R_CLK_posedge_posedge :	VitalDelayType := 2.200 ns;
      tsetup_S_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      thold_S_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      tpw_CLK_posedge :	VitalDelayType := 4.400 ns;
      tpw_R_negedge :	VitalDelayType := 4.400 ns;
      tperiod_CLK_posedge  :	VitalDelayType := 8.800 ns;
      ticd_CLK                       :	VitalDelayType := 0.000 ns;
      tisd_T_CLK                     :	VitalDelayType := 0.000 ns;
      tisd_R_CLK                     :	VitalDelayType := 0.000 ns;
      tisd_S_CLK                     :	VitalDelayType := 0.000 ns;
      tipd_T                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_R                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      T                              :	in    STD_ULOGIC;
      R                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of TFFRSS : entity is TRUE;
end TFFRSS;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library VF1;
architecture VITAL_VF of TFFRSS is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL T_ipd	 : STD_ULOGIC := 'X';
   SIGNAL R_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL T_CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL R_CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL S_CLK_dly	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (T_ipd, T, tipd_T);
   VitalWireDelay (R_ipd, R, tipd_R);
   VitalWireDelay (S_ipd, S, tipd_S);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   VitalSignalDelay (CLK_dly, CLK_ipd, ticd_CLK);
   VitalSignalDelay (T_CLK_dly, T_ipd, tisd_T_CLK);
   VitalSignalDelay (R_CLK_dly, R_ipd, tisd_R_CLK);
   VitalSignalDelay (S_CLK_dly, S_ipd, tisd_S_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (CLK_dly, T_CLK_dly, R_CLK_dly, S_CLK_dly)

   -- timing check results
   VARIABLE Tviol_T_CLK_R_EQ_1_ANB_S_EQ_1_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_T_CLK_R_EQ_1_ANB_S_EQ_1_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_R_CLK_S_EQ_1_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_R_CLK_S_EQ_1_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S_CLK_R_EQ_1_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S_CLK_R_EQ_1_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK_R_EQ_1_ANB_S_EQ_1	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK_R_EQ_1_ANB_S_EQ_1	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_R     : STD_ULOGIC := '0';
   VARIABLE PInfo_R     : VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 3);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;
   VARIABLE NOT_S_zd : STD_ULOGIC := '0';
   VARIABLE T_in_zd : STD_ULOGIC := '0';
   VARIABLE D_in_zd : STD_ULOGIC := '0';

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_T_CLK_R_EQ_1_ANB_S_EQ_1_posedge,
          TimingData              => Tmkr_T_CLK_R_EQ_1_ANB_S_EQ_1_posedge,
          TestSignal              => T_CLK_dly,
          TestSignalName          => "T",
          TestDelay               => tisd_T_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          SetupHigh               => tsetup_T_CLK_noedge_posedge,
          SetupLow                => tsetup_T_CLK_noedge_posedge,
          HoldHigh                => thold_T_CLK_noedge_posedge,
          HoldLow                 => thold_T_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((S_CLK_dly) AND (R_CLK_dly)) = '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/TFFRSS",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_R_CLK_S_EQ_1_posedge,
          TimingData              => Tmkr_R_CLK_S_EQ_1_posedge,
          TestSignal              => R_CLK_dly,
          TestSignalName          => "R",
          TestDelay               => tisd_R_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          Recovery                => trecovery_R_CLK_posedge_posedge,
          Removal                 => thold_R_CLK_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TO_X01(S_CLK_dly) = '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/TFFRSS",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_S_CLK_R_EQ_1_posedge,
          TimingData              => Tmkr_S_CLK_R_EQ_1_posedge,
          TestSignal              => S_CLK_dly,
          TestSignalName          => "S",
          TestDelay               => tisd_S_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          SetupHigh               => tsetup_S_CLK_noedge_posedge,
          SetupLow                => tsetup_S_CLK_noedge_posedge,
          HoldHigh                => thold_S_CLK_noedge_posedge,
          HoldLow                 => thold_S_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(R_CLK_dly) = '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/TFFRSS",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_R,
          PeriodData              => PInfo_R,
          TestSignal              => R_CLK_dly,
          TestSignalName          => "R",
          TestDelay               => tisd_R_CLK,
          Period                  => 0 ns,
          PulseWidthHigh          => tpw_R_negedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => TRUE,
          HeaderMsg               => InstancePath & "/TFFRSS",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK_R_EQ_1_ANB_S_EQ_1,
          PeriodData              => PInfo_CLK_R_EQ_1_ANB_S_EQ_1,
          TestSignal              => CLK_dly,
          TestSignalName          => "CLK",
          TestDelay               => ticd_CLK,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TO_X01(( (S_CLK_dly) ) AND ( (R_CLK_dly) )) = '1',
          HeaderMsg               => InstancePath & "/TFFRSS",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
        NOT_S_zd := VitalINV (S_CLK_dly);
        T_in_zd := VitalXOR2 (Q_zd, T_CLK_dly);
        D_in_zd := VitalOR2 (NOT_S_zd, T_in_zd);

      Violation := Tviol_T_CLK_R_EQ_1_ANB_S_EQ_1_posedge or Tviol_R_CLK_S_EQ_1_posedge or Tviol_S_CLK_R_EQ_1_posedge or Pviol_CLK_R_EQ_1_ANB_S_EQ_1;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => dfftab,
        DataIn => (
               D_in_zd, CLK_dly, R_CLK_dly, '1'));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (S_CLK_dly'last_event, tpd_S_Q, TRUE),
                 1 => (R_CLK_dly'last_event, tpd_R_Q, TRUE),
                 2 => (CLK_dly'last_event, tpd_CLK_Q, TRUE)),
       Mode => VitalInertial,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;

configuration CFG_TFFRSS_VITAL of TFFRSS is 
        for VITAL_VF
        end for; 
end CFG_TFFRSS_VITAL;
----- VITAL model for cell TFFRSSH -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;

LIBRARY VF1 ;
use VF1.VLOGTOVITAL_TABLES.all;



-- entity declaration --
entity TFFRSSH is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_S_Q                        :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tpd_R_Q                        :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tsetup_T_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      thold_T_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      trecovery_R_CLK_negedge_posedge :	VitalDelayType := 2.200 ns;
      thold_R_CLK_negedge_posedge :	VitalDelayType := 2.200 ns;
      tsetup_S_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      thold_S_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      tpw_CLK_posedge :	VitalDelayType := 4.400 ns;
      tpw_R_posedge :	VitalDelayType := 4.400 ns;
      tperiod_CLK_posedge  :	VitalDelayType := 8.800 ns;
      ticd_CLK                       :	VitalDelayType := 0.000 ns;
      tisd_T_CLK                     :	VitalDelayType := 0.000 ns;
      tisd_R_CLK                     :	VitalDelayType := 0.000 ns;
      tisd_S_CLK                     :	VitalDelayType := 0.000 ns;
      tipd_T                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_R                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      T                              :	in    STD_ULOGIC;
      R                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of TFFRSSH : entity is TRUE;
end TFFRSSH;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library VF1;
architecture VITAL_VF of TFFRSSH is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL T_ipd	 : STD_ULOGIC := 'X';
   SIGNAL R_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL T_CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL R_CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL S_CLK_dly	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (T_ipd, T, tipd_T);
   VitalWireDelay (R_ipd, R, tipd_R);
   VitalWireDelay (S_ipd, S, tipd_S);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   VitalSignalDelay (CLK_dly, CLK_ipd, ticd_CLK);
   VitalSignalDelay (T_CLK_dly, T_ipd, tisd_T_CLK);
   VitalSignalDelay (R_CLK_dly, R_ipd, tisd_R_CLK);
   VitalSignalDelay (S_CLK_dly, S_ipd, tisd_S_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (CLK_dly, T_CLK_dly, R_CLK_dly, S_CLK_dly)

   -- timing check results
   VARIABLE Tviol_T_CLK_R_EQ_0_ANB_S_EQ_0_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_T_CLK_R_EQ_0_ANB_S_EQ_0_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_R_CLK_S_EQ_0_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_R_CLK_S_EQ_0_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S_CLK_R_EQ_0_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S_CLK_R_EQ_0_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK_R_EQ_0_ANB_S_EQ_0	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK_R_EQ_0_ANB_S_EQ_0	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_R     : STD_ULOGIC := '0';
   VARIABLE PInfo_R     : VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 3);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');

   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;
   VARIABLE NOT_S_zd : STD_ULOGIC := '0';
   VARIABLE R_inverted : STD_ULOGIC := 'X';
   VARIABLE T_in_zd : STD_ULOGIC := '0';
   VARIABLE D_in_zd : STD_ULOGIC := '0';

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_T_CLK_R_EQ_0_ANB_S_EQ_0_posedge,
          TimingData              => Tmkr_T_CLK_R_EQ_0_ANB_S_EQ_0_posedge,
          TestSignal              => T_CLK_dly,
          TestSignalName          => "T",
          TestDelay               => tisd_T_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          SetupHigh               => tsetup_T_CLK_noedge_posedge,
          SetupLow                => tsetup_T_CLK_noedge_posedge,
          HoldHigh                => thold_T_CLK_noedge_posedge,
          HoldLow                 => thold_T_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(((NOT S_CLK_dly)) AND ((NOT R_CLK_dly))) = '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/TFFRSSH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_R_CLK_S_EQ_0_posedge,
          TimingData              => Tmkr_R_CLK_S_EQ_0_posedge,
          TestSignal              => R_CLK_dly,
          TestSignalName          => "R",
          TestDelay               => tisd_R_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          Recovery                => trecovery_R_CLK_negedge_posedge,
          Removal                 => thold_R_CLK_negedge_posedge,
          ActiveLow               => FALSE,
          CheckEnabled            => 
                           TO_X01((S_CLK_dly)) = '0',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/TFFRSSH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_S_CLK_R_EQ_0_posedge,
          TimingData              => Tmkr_S_CLK_R_EQ_0_posedge,
          TestSignal              => S_CLK_dly,
          TestSignalName          => "S",
          TestDelay               => tisd_S_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          SetupHigh               => tsetup_S_CLK_noedge_posedge,
          SetupLow                => tsetup_S_CLK_noedge_posedge,
          HoldHigh                => thold_S_CLK_noedge_posedge,
          HoldLow                 => thold_S_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((R_CLK_dly)) = '0',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/TFFRSSH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_R,
          PeriodData              => PInfo_R,
          TestSignal              => R_CLK_dly,
          TestSignalName          => "R",
          TestDelay               => tisd_R_CLK,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_R_posedge,
          CheckEnabled            => TRUE, 
          HeaderMsg               => InstancePath & "/TFFRSSH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK_R_EQ_0_ANB_S_EQ_0,
          PeriodData              => PInfo_CLK_R_EQ_0_ANB_S_EQ_0,
          TestSignal              => CLK_dly,
          TestSignalName          => "CLK",
          TestDelay               => ticd_CLK,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TO_X01(( NOT S_CLK_dly ) AND ( NOT R_CLK_dly ) ) = '1',
          HeaderMsg               => InstancePath & "/TFFRSSH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
        R_inverted := NOT (R_CLK_dly);
        T_in_zd := VitalXOR2 (Q_zd, T_CLK_dly);
        D_in_zd := VitalOR2 (S_CLK_dly, T_in_zd);

      Violation := Tviol_T_CLK_R_EQ_0_ANB_S_EQ_0_posedge or Tviol_R_CLK_S_EQ_0_posedge or Tviol_S_CLK_R_EQ_0_posedge or Pviol_CLK_R_EQ_0_ANB_S_EQ_0 or Pviol_R;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => dfftab,
        DataIn => (
               D_in_zd, CLK_dly, R_inverted, '1'));
        Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (S_CLK_dly'last_event, tpd_S_Q, TRUE),
                 1 => (R_CLK_dly'last_event, tpd_R_Q, TRUE),
                 2 => (CLK_dly'last_event, tpd_CLK_Q, TRUE)),
       Mode => VitalInertial,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;

configuration CFG_TFFRSSH_VITAL of TFFRSSH is 
        for VITAL_VF
        end for; 
end CFG_TFFRSSH_VITAL;
----- VITAL model for cell TFFS -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;

LIBRARY VF1 ;
use VF1.VLOGTOVITAL_TABLES.all;



-- entity declaration --
entity TFFS is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_S_Q                        :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tsetup_T_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      thold_T_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      trecovery_S_CLK_posedge_posedge :	VitalDelayType := 2.200 ns;
      thold_S_CLK_posedge_posedge    :	VitalDelayType := 2.200 ns;
      tpw_CLK_posedge         :	VitalDelayType := 4.400 ns;
      tperiod_CLK_posedge             :	VitalDelayType := 8.800 ns;
      ticd_CLK                       :	VitalDelayType := 0.000 ns;
      tisd_T_CLK                     :	VitalDelayType := 0.000 ns;
      tisd_S_CLK                     :	VitalDelayType := 0.000 ns;
      tipd_T                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      T                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of TFFS : entity is TRUE;
end TFFS;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library VF1;
architecture VITAL_VF of TFFS is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL T_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL T_CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL S_CLK_dly	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (T_ipd, T, tipd_T);
   VitalWireDelay (S_ipd, S, tipd_S);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   VitalSignalDelay (CLK_dly, CLK_ipd, ticd_CLK);
   VitalSignalDelay (T_CLK_dly, T_ipd, tisd_T_CLK);
   VitalSignalDelay (S_CLK_dly, S_ipd, tisd_S_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (CLK_dly, T_CLK_dly, S_CLK_dly)

   -- timing check results
   VARIABLE Tviol_T_CLK_S_EQ_1_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_T_CLK_S_EQ_1_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK_S_EQ_1	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK_S_EQ_1	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 3);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_T_CLK_S_EQ_1_posedge,
          TimingData              => Tmkr_T_CLK_S_EQ_1_posedge,
          TestSignal              => T_CLK_dly,
          TestSignalName          => "T",
          TestDelay               => tisd_T_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          SetupHigh               => tsetup_T_CLK_noedge_posedge,
          SetupLow                => tsetup_T_CLK_noedge_posedge,
          HoldHigh                => thold_T_CLK_noedge_posedge,
          HoldLow                 => thold_T_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(S_CLK_dly) = '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/TFFS",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_S_CLK_posedge,
          TimingData              => Tmkr_S_CLK_posedge,
          TestSignal              => S_CLK_dly,
          TestSignalName          => "S",
          TestDelay               => tisd_S_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          Recovery                => trecovery_S_CLK_posedge_posedge,
          Removal                 => thold_S_CLK_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/TFFS",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK_S_EQ_1,
          PeriodData              => PInfo_CLK_S_EQ_1,
          TestSignal              => CLK_dly,
          TestSignalName          => "CLK",
          TestDelay               => ticd_CLK,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TO_X01((S_CLK_dly) ) = '1',
          HeaderMsg               => InstancePath & "/TFFS",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_T_CLK_S_EQ_1_posedge or Tviol_S_CLK_posedge or Pviol_CLK_S_EQ_1;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => tfftab,
        DataIn => (
               CLK_dly, T_CLK_dly, S_CLK_dly, '1'));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (S_CLK_dly'last_event, tpd_S_Q, TRUE),
                 1 => (CLK_dly'last_event, tpd_CLK_Q, TRUE)),
       Mode => VitalInertial,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;

configuration CFG_TFFS_VITAL of TFFS is 
        for VITAL_VF
        end for; 
end CFG_TFFS_VITAL;
----- VITAL model for cell TFFSH -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;

LIBRARY VF1 ;
use VF1.VLOGTOVITAL_TABLES.all;



-- entity declaration --
entity TFFSH is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_S_Q                        :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.440 ns, 1.440 ns);
      tsetup_T_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      thold_T_CLK_noedge_posedge :	VitalDelayType := 2.200 ns;
      trecovery_S_CLK_negedge_posedge :	VitalDelayType := 2.200 ns;
      thold_S_CLK_negedge_posedge    :	VitalDelayType := 2.200 ns;
      tpw_CLK_posedge         :	VitalDelayType := 4.400 ns;
      tpw_S_posedge         :	VitalDelayType := 4.400 ns;
      tperiod_CLK_posedge             :	VitalDelayType := 8.800 ns;
      ticd_CLK                       :	VitalDelayType := 0.000 ns;
      tisd_T_CLK                     :	VitalDelayType := 0.000 ns;
      tisd_S_CLK                     :	VitalDelayType := 0.000 ns;
      tipd_T                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      T                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of TFFSH : entity is TRUE;
end TFFSH;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library VF1;
architecture VITAL_VF of TFFSH is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL T_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL T_CLK_dly	 : STD_ULOGIC := 'X';
   SIGNAL S_CLK_dly	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (T_ipd, T, tipd_T);
   VitalWireDelay (S_ipd, S, tipd_S);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   VitalSignalDelay (CLK_dly, CLK_ipd, ticd_CLK);
   VitalSignalDelay (T_CLK_dly, T_ipd, tisd_T_CLK);
   VitalSignalDelay (S_CLK_dly, S_ipd, tisd_S_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (CLK_dly, T_CLK_dly, S_CLK_dly)

   -- timing check results
   VARIABLE Tviol_T_CLK_S_EQ_0_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_T_CLK_S_EQ_0_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK_S_EQ_0	: STD_ULOGIC := '0';
   VARIABLE Pviol_S	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK_S_EQ_0	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE PInfo_S	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 3);
   VARIABLE S_inverted : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_T_CLK_S_EQ_0_posedge,
          TimingData              => Tmkr_T_CLK_S_EQ_0_posedge,
          TestSignal              => T_CLK_dly,
          TestSignalName          => "T",
          TestDelay               => tisd_T_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          SetupHigh               => tsetup_T_CLK_noedge_posedge,
          SetupLow                => tsetup_T_CLK_noedge_posedge,
          HoldHigh                => thold_T_CLK_noedge_posedge,
          HoldLow                 => thold_T_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((S_CLK_dly)) = '0',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/TFFSH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_S_CLK_posedge,
          TimingData              => Tmkr_S_CLK_posedge,
          TestSignal              => S_CLK_dly,
          TestSignalName          => "S",
          TestDelay               => tisd_S_CLK,
          RefSignal               => CLK_dly,
          RefSignalName          => "CLK",
          RefDelay                => ticd_CLK,
          Recovery                => trecovery_S_CLK_negedge_posedge,
          Removal                 => thold_S_CLK_negedge_posedge,
          ActiveLow               => FALSE,
          CheckEnabled            => TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/TFFSH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_S,
          PeriodData              => PInfo_S,
          TestSignal              => S_CLK_dly,
          TestSignalName          => "S",
          TestDelay               => tisd_S_CLK,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_S_posedge,
          CheckEnabled            => TRUE, 
          HeaderMsg               => InstancePath & "/TFFSH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK_S_EQ_0,
          PeriodData              => PInfo_CLK_S_EQ_0,
          TestSignal              => CLK_dly,
          TestSignalName          => "CLK",
          TestDelay               => ticd_CLK,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TO_X01(S_CLK_dly ) = '0',
          HeaderMsg               => InstancePath & "/TFFSH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_T_CLK_S_EQ_0_posedge or Tviol_S_CLK_posedge or Pviol_CLK_S_EQ_0 or Pviol_S;
      S_inverted := (NOT S_CLK_dly);
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => tfftab,
        DataIn => (
               CLK_dly, T_CLK_dly, S_inverted, '1'));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (S_CLK_dly'last_event, tpd_S_Q, TRUE),
                 1 => (CLK_dly'last_event, tpd_CLK_Q, TRUE)),
       Mode => VitalInertial,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;

configuration CFG_TFFSH_VITAL of TFFSH is 
        for VITAL_VF
        end for; 
end CFG_TFFSH_VITAL;
----- VITAL model for cell VCC -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity VCC is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True);

   port(
      X                              :	out   STD_ULOGIC := '1');
attribute VITAL_LEVEL0 of VCC : entity is TRUE;
end VCC;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library VF1;
architecture VITAL_VF of VCC is
   attribute VITAL_LEVEL0 of VITAL_VF : architecture is TRUE;
   
   SIGNAL SUPPLY1  : STD_ULOGIC := '1'; 

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   --  empty
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------

Inst1: VitalBUF (X,SUPPLY1);

end VITAL_VF;

configuration CFG_VCC_VITAL of VCC is 
        for VITAL_VF
        end for; 
end CFG_VCC_VITAL;
----- VITAL model for cell XNOR2 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity XNOR2 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_I0_O                       :	VitalDelayType01 := (1.25 ns, 1.25 ns);
      tpd_I1_O                       :	VitalDelayType01 := (1.25 ns, 1.25 ns);
      tipd_I0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      I0                             :	in    STD_ULOGIC;
      I1                             :	in    STD_ULOGIC;
      O                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of XNOR2 : entity is TRUE;
end XNOR2;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library VF1;
architecture VITAL_VF of XNOR2 is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL I0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I1_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (I0_ipd, I0, tipd_I0);
   VitalWireDelay (I1_ipd, I1, tipd_I1);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (I0_ipd, I1_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS O_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE O_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      O_zd :=
       (((NOT I1_ipd)) AND ((NOT I0_ipd))) OR ((I1_ipd) AND (I0_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => O,
       GlitchData => O_GlitchData,
       OutSignalName => "O",
       OutTemp => O_zd,
       Paths => (0 => (I0_ipd'last_event, tpd_I0_O, TRUE),
                 1 => (I1_ipd'last_event, tpd_I1_O, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;

configuration CFG_XNOR2_VITAL of XNOR2 is 
        for VITAL_VF
        end for; 
end CFG_XNOR2_VITAL;
----- VITAL model for cell XNOR3 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity XNOR3 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_I0_O                       :	VitalDelayType01 := (1.250 ns, 1.250 ns);
      tpd_I1_O                       :	VitalDelayType01 := (1.250 ns, 1.250 ns);
      tpd_I2_O                       :	VitalDelayType01 := (1.250 ns, 1.250 ns);
      tipd_I0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I2                        :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      I0                             :	in    STD_ULOGIC;
      I1                             :	in    STD_ULOGIC;
      I2                             :	in    STD_ULOGIC;
      O                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of XNOR3 : entity is TRUE;
end XNOR3;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_VF of XNOR3 is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL I0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I1_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I2_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (I0_ipd, I0, tipd_I0);
   VitalWireDelay (I1_ipd, I1, tipd_I1);
   VitalWireDelay (I2_ipd, I2, tipd_I2);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (I0_ipd, I1_ipd, I2_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS O_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE O_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      O_zd := (NOT ((I1_ipd) XOR (I0_ipd) XOR (I2_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => O,
       GlitchData => O_GlitchData,
       OutSignalName => "O",
       OutTemp => O_zd,
       Paths => (0 => (I0_ipd'last_event, tpd_I0_O, TRUE),
                 1 => (I1_ipd'last_event, tpd_I1_O, TRUE),
                 2 => (I2_ipd'last_event, tpd_I2_O, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;

configuration CFG_XNOR3_VITAL of XNOR3 is 
        for VITAL_VF
        end for; 
end CFG_XNOR3_VITAL;
----- VITAL model for cell XNOR4 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity XNOR4 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_I0_O                       :	VitalDelayType01 := (1.800 ns, 1.800 ns);
      tpd_I1_O                       :	VitalDelayType01 := (1.800 ns, 1.800 ns);
      tpd_I2_O                       :	VitalDelayType01 := (1.800 ns, 1.800 ns);
      tpd_I3_O                       :	VitalDelayType01 := (1.800 ns, 1.800 ns);
      tipd_I0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I2                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I3                        :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      I0                             :	in    STD_ULOGIC;
      I1                             :	in    STD_ULOGIC;
      I2                             :	in    STD_ULOGIC;
      I3                             :	in    STD_ULOGIC;
      O                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of XNOR4 : entity is TRUE;
end XNOR4;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_VF of XNOR4 is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL I0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I1_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I2_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I3_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (I0_ipd, I0, tipd_I0);
   VitalWireDelay (I1_ipd, I1, tipd_I1);
   VitalWireDelay (I2_ipd, I2, tipd_I2);
   VitalWireDelay (I3_ipd, I3, tipd_I3);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (I0_ipd, I1_ipd, I2_ipd, I3_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS O_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE O_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      O_zd := (NOT ((I1_ipd) XOR (I0_ipd) XOR (I2_ipd) XOR (I3_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => O,
       GlitchData => O_GlitchData,
       OutSignalName => "O",
       OutTemp => O_zd,
       Paths => (0 => (I0_ipd'last_event, tpd_I0_O, TRUE),
                 1 => (I1_ipd'last_event, tpd_I1_O, TRUE),
                 2 => (I2_ipd'last_event, tpd_I2_O, TRUE),
                 3 => (I3_ipd'last_event, tpd_I3_O, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;

configuration CFG_XNOR4_VITAL of XNOR4 is 
        for VITAL_VF
        end for; 
end CFG_XNOR4_VITAL;
----- VITAL model for cell XNOR5 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity XNOR5 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_I0_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I1_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I2_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I3_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I4_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tipd_I0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I2                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I3                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I4                        :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      I0                             :	in    STD_ULOGIC;
      I1                             :	in    STD_ULOGIC;
      I2                             :	in    STD_ULOGIC;
      I3                             :	in    STD_ULOGIC;
      I4                             :	in    STD_ULOGIC;
      O                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of XNOR5 : entity is TRUE;
end XNOR5;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
 
library VF1;
architecture VITAL_VF of XNOR5 is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL I0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I1_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I2_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I3_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I4_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (I0_ipd, I0, tipd_I0);
   VitalWireDelay (I1_ipd, I1, tipd_I1);
   VitalWireDelay (I2_ipd, I2, tipd_I2);
   VitalWireDelay (I3_ipd, I3, tipd_I3);
   VitalWireDelay (I4_ipd, I4, tipd_I4);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (I0_ipd, I1_ipd, I2_ipd, I3_ipd, I4_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS O_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE O_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      O_zd :=
       (NOT ((I1_ipd) XOR (I0_ipd) XOR (I2_ipd) XOR (I3_ipd) XOR (I4_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => O,
       GlitchData => O_GlitchData,
       OutSignalName => "O",
       OutTemp => O_zd,
       Paths => (0 => (I0_ipd'last_event, tpd_I0_O, TRUE),
                 1 => (I1_ipd'last_event, tpd_I1_O, TRUE),
                 2 => (I2_ipd'last_event, tpd_I2_O, TRUE),
                 3 => (I3_ipd'last_event, tpd_I3_O, TRUE),
                 4 => (I4_ipd'last_event, tpd_I4_O, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;
 
configuration CFG_XNOR5_VITAL of XNOR5 is 
        for VITAL_VF
        end for; 
end CFG_XNOR5_VITAL;
----- VITAL model for cell XNOR6 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity XNOR6 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_I0_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I1_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I2_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I3_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I4_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I5_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tipd_I0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I2                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I3                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I4                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I5                        :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      I0                             :	in    STD_ULOGIC;
      I1                             :	in    STD_ULOGIC;
      I2                             :	in    STD_ULOGIC;
      I3                             :	in    STD_ULOGIC;
      I4                             :	in    STD_ULOGIC;
      I5                             :	in    STD_ULOGIC;
      O                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of XNOR6 : entity is TRUE;
end XNOR6;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
 
library VF1;
architecture VITAL_VF of XNOR6 is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL I0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I1_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I2_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I3_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I4_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I5_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (I0_ipd, I0, tipd_I0);
   VitalWireDelay (I1_ipd, I1, tipd_I1);
   VitalWireDelay (I2_ipd, I2, tipd_I2);
   VitalWireDelay (I3_ipd, I3, tipd_I3);
   VitalWireDelay (I4_ipd, I4, tipd_I4);
   VitalWireDelay (I5_ipd, I5, tipd_I5);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (I0_ipd, I1_ipd, I2_ipd, I3_ipd, I4_ipd, I5_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS O_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE O_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      O_zd :=
       (NOT ((I1_ipd) XOR (I0_ipd) XOR (I2_ipd) XOR (I3_ipd) XOR (I4_ipd)
         XOR (I5_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => O,
       GlitchData => O_GlitchData,
       OutSignalName => "O",
       OutTemp => O_zd,
       Paths => (0 => (I0_ipd'last_event, tpd_I0_O, TRUE),
                 1 => (I1_ipd'last_event, tpd_I1_O, TRUE),
                 2 => (I2_ipd'last_event, tpd_I2_O, TRUE),
                 3 => (I3_ipd'last_event, tpd_I3_O, TRUE),
                 4 => (I4_ipd'last_event, tpd_I4_O, TRUE),
                 5 => (I5_ipd'last_event, tpd_I5_O, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;
 
configuration CFG_XNOR6_VITAL of XNOR6 is 
        for VITAL_VF
        end for; 
end CFG_XNOR6_VITAL;
----- VITAL model for cell XOR2 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity XOR2 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_I0_O                       :	VitalDelayType01 := (1.25 ns, 1.25 ns);
      tpd_I1_O                       :	VitalDelayType01 := (1.25 ns, 1.25 ns);
      tipd_I0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      I0                             :	in    STD_ULOGIC;
      I1                             :	in    STD_ULOGIC;
      O                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of XOR2 : entity is TRUE;

   -- real names
   -- REAL_NAME of XOR2 is "XOR2"
end XOR2;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library VF1;
architecture VITAL_VF of XOR2 is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL I0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I1_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (I0_ipd, I0, tipd_I0);
   VitalWireDelay (I1_ipd, I1, tipd_I1);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (I0_ipd, I1_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS O_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE O_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      O_zd :=
       (((NOT I0_ipd)) AND (I1_ipd)) OR (((NOT I1_ipd)) AND (I0_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => O,
       GlitchData => O_GlitchData,
       OutSignalName => "O",
       OutTemp => O_zd,
       Paths => (0 => (I0_ipd'last_event, tpd_I0_O, TRUE),
                 1 => (I1_ipd'last_event, tpd_I1_O, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;

configuration CFG_XOR2_VITAL of XOR2 is 
        for VITAL_VF
        end for; 
end CFG_XOR2_VITAL;
----- VITAL model for cell XOR3 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity XOR3 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_I0_O                       :	VitalDelayType01 := (1.250 ns, 1.250 ns);
      tpd_I1_O                       :	VitalDelayType01 := (1.250 ns, 1.250 ns);
      tpd_I2_O                       :	VitalDelayType01 := (1.250 ns, 1.250 ns);
      tipd_I0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I2                        :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      I0                             :	in    STD_ULOGIC;
      I1                             :	in    STD_ULOGIC;
      I2                             :	in    STD_ULOGIC;
      O                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of XOR3 : entity is TRUE;
end XOR3;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_VF of XOR3 is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL I0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I1_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I2_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (I0_ipd, I0, tipd_I0);
   VitalWireDelay (I1_ipd, I1, tipd_I1);
   VitalWireDelay (I2_ipd, I2, tipd_I2);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (I0_ipd, I1_ipd, I2_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS O_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE O_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      O_zd := (I1_ipd) XOR (I0_ipd) XOR (I2_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => O,
       GlitchData => O_GlitchData,
       OutSignalName => "O",
       OutTemp => O_zd,
       Paths => (0 => (I0_ipd'last_event, tpd_I0_O, TRUE),
                 1 => (I1_ipd'last_event, tpd_I1_O, TRUE),
                 2 => (I2_ipd'last_event, tpd_I2_O, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;

configuration CFG_XOR3_VITAL of XOR3 is 
        for VITAL_VF
        end for; 
end CFG_XOR3_VITAL;
----- VITAL model for cell XOR4 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity XOR4 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_I0_O                       :	VitalDelayType01 := (1.800 ns, 1.800 ns);
      tpd_I1_O                       :	VitalDelayType01 := (1.800 ns, 1.800 ns);
      tpd_I2_O                       :	VitalDelayType01 := (1.800 ns, 1.800 ns);
      tpd_I3_O                       :	VitalDelayType01 := (1.800 ns, 1.800 ns);
      tipd_I0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I2                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I3                        :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      I0                             :	in    STD_ULOGIC;
      I1                             :	in    STD_ULOGIC;
      I2                             :	in    STD_ULOGIC;
      I3                             :	in    STD_ULOGIC;
      O                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of XOR4 : entity is TRUE;
end XOR4;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_VF of XOR4 is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL I0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I1_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I2_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I3_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (I0_ipd, I0, tipd_I0);
   VitalWireDelay (I1_ipd, I1, tipd_I1);
   VitalWireDelay (I2_ipd, I2, tipd_I2);
   VitalWireDelay (I3_ipd, I3, tipd_I3);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (I0_ipd, I1_ipd, I2_ipd, I3_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS O_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE O_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      O_zd := (I1_ipd) XOR (I0_ipd) XOR (I2_ipd) XOR (I3_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => O,
       GlitchData => O_GlitchData,
       OutSignalName => "O",
       OutTemp => O_zd,
       Paths => (0 => (I0_ipd'last_event, tpd_I0_O, TRUE),
                 1 => (I1_ipd'last_event, tpd_I1_O, TRUE),
                 2 => (I2_ipd'last_event, tpd_I2_O, TRUE),
                 3 => (I3_ipd'last_event, tpd_I3_O, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;

configuration CFG_XOR4_VITAL of XOR4 is 
        for VITAL_VF
        end for; 
end CFG_XOR4_VITAL;
----- VITAL model for cell XOR5 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity XOR5 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_I0_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I1_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I2_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I3_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I4_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tipd_I0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I2                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I3                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I4                        :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      I0                             :	in    STD_ULOGIC;
      I1                             :	in    STD_ULOGIC;
      I2                             :	in    STD_ULOGIC;
      I3                             :	in    STD_ULOGIC;
      I4                             :	in    STD_ULOGIC;
      O                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of XOR5 : entity is TRUE;
end XOR5;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
 
library VF1;
architecture VITAL_VF of XOR5 is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL I0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I1_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I2_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I3_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I4_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (I0_ipd, I0, tipd_I0);
   VitalWireDelay (I1_ipd, I1, tipd_I1);
   VitalWireDelay (I2_ipd, I2, tipd_I2);
   VitalWireDelay (I3_ipd, I3, tipd_I3);
   VitalWireDelay (I4_ipd, I4, tipd_I4);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (I0_ipd, I1_ipd, I2_ipd, I3_ipd, I4_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS O_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE O_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      O_zd :=
       (I1_ipd) XOR (I0_ipd) XOR (I2_ipd) XOR (I3_ipd) XOR (I4_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => O,
       GlitchData => O_GlitchData,
       OutSignalName => "O",
       OutTemp => O_zd,
       Paths => (0 => (I0_ipd'last_event, tpd_I0_O, TRUE),
                 1 => (I1_ipd'last_event, tpd_I1_O, TRUE),
                 2 => (I2_ipd'last_event, tpd_I2_O, TRUE),
                 3 => (I3_ipd'last_event, tpd_I3_O, TRUE),
                 4 => (I4_ipd'last_event, tpd_I4_O, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;
 
configuration CFG_XOR5_VITAL of XOR5 is 
        for VITAL_VF
        end for; 
end CFG_XOR5_VITAL;
----- VITAL model for cell XOR6 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity XOR6 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_I0_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I1_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I2_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I3_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I4_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tpd_I5_O                       :	VitalDelayType01 := (2.500 ns, 2.500 ns);
      tipd_I0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I2                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I3                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I4                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I5                        :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      I0                             :	in    STD_ULOGIC;
      I1                             :	in    STD_ULOGIC;
      I2                             :	in    STD_ULOGIC;
      I3                             :	in    STD_ULOGIC;
      I4                             :	in    STD_ULOGIC;
      I5                             :	in    STD_ULOGIC;
      O                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of XOR6 : entity is TRUE;
end XOR6;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
 
library VF1;
architecture VITAL_VF of XOR6 is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL I0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I1_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I2_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I3_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I4_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I5_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (I0_ipd, I0, tipd_I0);
   VitalWireDelay (I1_ipd, I1, tipd_I1);
   VitalWireDelay (I2_ipd, I2, tipd_I2);
   VitalWireDelay (I3_ipd, I3, tipd_I3);
   VitalWireDelay (I4_ipd, I4, tipd_I4);
   VitalWireDelay (I5_ipd, I5, tipd_I5);
   end block;
   ----------------------
   --  INPUT SIGNAL DELAYs
   ----------------------
   SignalDelay : block
   begin
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (I0_ipd, I1_ipd, I2_ipd, I3_ipd, I4_ipd, I5_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS O_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE O_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      O_zd :=
       (I1_ipd) XOR (I0_ipd) XOR (I2_ipd) XOR (I3_ipd) XOR (I4_ipd) XOR
         (I5_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => O,
       GlitchData => O_GlitchData,
       OutSignalName => "O",
       OutTemp => O_zd,
       Paths => (0 => (I0_ipd'last_event, tpd_I0_O, TRUE),
                 1 => (I1_ipd'last_event, tpd_I1_O, TRUE),
                 2 => (I2_ipd'last_event, tpd_I2_O, TRUE),
                 3 => (I3_ipd'last_event, tpd_I3_O, TRUE),
                 4 => (I4_ipd'last_event, tpd_I4_O, TRUE),
                 5 => (I5_ipd'last_event, tpd_I5_O, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;
 
configuration CFG_XOR6_VITAL of XOR6 is 
        for VITAL_VF
        end for; 
end CFG_XOR6_VITAL;
----- VITAL model for cell XORSOFT -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity XORSOFT is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_I0_O                       :	VitalDelayType01 := (1.25 ns, 1.25 ns);
      tpd_I1_O                       :	VitalDelayType01 := (1.25 ns, 1.25 ns);
      tipd_I0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_I1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      I0                             :	in    STD_ULOGIC;
      I1                             :	in    STD_ULOGIC;
      O                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of XORSOFT : entity is TRUE;
end XORSOFT;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library VF1;
architecture VITAL_VF of XORSOFT is
   attribute VITAL_LEVEL1 of VITAL_VF : architecture is TRUE;

   SIGNAL I0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL I1_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (I0_ipd, I0, tipd_I0);
   VitalWireDelay (I1_ipd, I1, tipd_I1);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (I0_ipd, I1_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS O_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE O_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      O_zd :=
       (((NOT I0_ipd)) AND (I1_ipd)) OR (((NOT I1_ipd)) AND (I0_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => O,
       GlitchData => O_GlitchData,
       OutSignalName => "O",
       OutTemp => O_zd,
       Paths => (0 => (I0_ipd'last_event, tpd_I0_O, TRUE),
                 1 => (I1_ipd'last_event, tpd_I1_O, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL_VF;

configuration CFG_XORSOFT_VITAL of XORSOFT is 
        for VITAL_VF
        end for; 
end CFG_XORSOFT_VITAL;
-----------------------------------------------------------------------
-- Local Package
-----------------------------------------------------------------------

LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
LIBRARY VF1;
USE VF1.ALL;

package RAMPACK is

  subtype data_word_typ is std_logic_vector (3 downto 0);
  subtype address_type is std_logic_vector (4 downto 0);
  type memory_array_typ is array(0 to 31) of data_word_typ;

  constant x_data : data_word_typ := ('X','X','X','X');
  constant z_data : data_word_typ := ('Z','Z','Z','Z');
  constant x_add : address_type := ('X','X','X','X','X');

   function vec2int		(v:	std_logic_vector)	return integer;

   function bitX		(v:	std_logic)		return boolean;

   function vecX		(v:	std_logic_vector)	return boolean;

end;

package body RAMPACK is

------------------------------------------------------------------------
   function vec2int           (v: std_logic_vector) return integer is
      variable result: integer := 0;
      variable addition: integer := 1;
   begin
      for b in v'reverse_range loop
         if v (b) = '1' then
            result := result + addition;
         end if;
         addition := addition * 2;
      end loop;
      return result;
   end;

------------------------------------------------------------------------

------------------------------------------------------------------------
   function vecX              (v:        std_logic_vector) return boolean is
   begin
      for b in v'range loop
         if bitX (v (b)) then
            return true;
         end if;
      end loop;
      return false;
   end;

------------------------------------------------------------------------

------------------------------------------------------------------------
   function bitX              (v:        std_logic)    return boolean is
   begin
      case v is
         when 'X'    => return true;
         when others => return false;
      end case;
   end;

------------------------------------------------------------------------

end RAMPACK;
-------------------------------------------------------------------------------


---------------------------------------------------------------------
-- VITAL model for RB_DA 30.10 technology
-----------------------------------------------------------------------

LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.VITAL_timing.all;
USE IEEE.std_logic_textio.all;
USE IEEE.VITAL_primitives.all;
LIBRARY std;
USE std.textio.all;
LIBRARY VF1;
USE VF1.ALL;
USE VF1.RAMPACK.ALL;

-----------------------------------------------------------------------
-- ENTITY declaration
-----------------------------------------------------------------------

ENTITY RB_DA IS
  GENERIC (
	tipd_WEN		: VitalDelayType01			:= (0.0 ns, 0.0 ns);
	tipd_REN		: VitalDelayType01			:= (0.0 ns, 0.0 ns);
	tipd_WRCLK		: VitalDelayType01			:= (0.0 ns, 0.0 ns);
	tipd_OE		: VitalDelayType01			:= (0.0 ns, 0.0 ns);
        tipd_WRDATA3            : VitalDelayType01      := (0.0 ns, 0.0 ns);
        tipd_WRDATA2            : VitalDelayType01      := (0.0 ns, 0.0 ns);
        tipd_WRDATA1            : VitalDelayType01      := (0.0 ns, 0.0 ns);
        tipd_WRDATA0            : VitalDelayType01      := (0.0 ns, 0.0 ns);
        tipd_WRAD4              : VitalDelayType01      := (0.0 ns, 0.0 ns);
        tipd_WRAD3              : VitalDelayType01      := (0.0 ns, 0.0 ns);
        tipd_WRAD2              : VitalDelayType01      := (0.0 ns, 0.0 ns);
        tipd_WRAD1              : VitalDelayType01      := (0.0 ns, 0.0 ns);
        tipd_WRAD0              : VitalDelayType01      := (0.0 ns, 0.0 ns);
        tipd_RAD4              : VitalDelayType01      := (0.0 ns, 0.0 ns);
        tipd_RAD3              : VitalDelayType01      := (0.0 ns, 0.0 ns);
        tipd_RAD2              : VitalDelayType01      := (0.0 ns, 0.0 ns);
        tipd_RAD1              : VitalDelayType01      := (0.0 ns, 0.0 ns);
        tipd_RAD0              : VitalDelayType01      := (0.0 ns, 0.0 ns);

tpd_WRAD4_WRDATA0         :VitalDelayType01Z := (2 ns,2 ns,2 ns,2 ns,2 ns,2 ns);
tpd_WRAD3_WRDATA0         :VitalDelayType01Z := (2 ns,2 ns,2 ns,2 ns,2 ns,2 ns);
tpd_WRAD2_WRDATA0         :VitalDelayType01Z := (2 ns,2 ns,2 ns,2 ns,2 ns,2 ns);
tpd_WRAD1_WRDATA0         :VitalDelayType01Z := (2 ns,2 ns,2 ns,2 ns,2 ns,2 ns);
tpd_WRAD0_WRDATA0         :VitalDelayType01Z := (2 ns,2 ns,2 ns,2 ns,2 ns,2 ns);
tpd_WRAD4_WRDATA1         :VitalDelayType01Z := (2 ns,2 ns,2 ns,2 ns,2 ns,2 ns);
tpd_WRAD3_WRDATA1         :VitalDelayType01Z := (2 ns,2 ns,2 ns,2 ns,2 ns,2 ns);
tpd_WRAD2_WRDATA1         :VitalDelayType01Z := (2 ns,2 ns,2 ns,2 ns,2 ns,2 ns);
tpd_WRAD1_WRDATA1         :VitalDelayType01Z := (2 ns,2 ns,2 ns,2 ns,2 ns,2 ns);
tpd_WRAD0_WRDATA1         :VitalDelayType01Z := (2 ns,2 ns,2 ns,2 ns,2 ns,2 ns);
tpd_WRAD4_WRDATA2         :VitalDelayType01Z := (2 ns,2 ns,2 ns,2 ns,2 ns,2 ns);
tpd_WRAD3_WRDATA2         :VitalDelayType01Z := (2 ns,2 ns,2 ns,2 ns,2 ns,2 ns);
tpd_WRAD2_WRDATA2         :VitalDelayType01Z := (2 ns,2 ns,2 ns,2 ns,2 ns,2 ns);
tpd_WRAD1_WRDATA2         :VitalDelayType01Z := (2 ns,2 ns,2 ns,2 ns,2 ns,2 ns);
tpd_WRAD0_WRDATA2         :VitalDelayType01Z := (2 ns,2 ns,2 ns,2 ns,2 ns,2 ns);
tpd_WRAD4_WRDATA3         :VitalDelayType01Z := (2 ns,2 ns,2 ns,2 ns,2 ns,2 ns);
tpd_WRAD3_WRDATA3         :VitalDelayType01Z := (2 ns,2 ns,2 ns,2 ns,2 ns,2 ns);
tpd_WRAD2_WRDATA3         :VitalDelayType01Z := (2 ns,2 ns,2 ns,2 ns,2 ns,2 ns);
tpd_WRAD1_WRDATA3         :VitalDelayType01Z := (2 ns,2 ns,2 ns,2 ns,2 ns,2 ns);
tpd_WRAD0_WRDATA3         :VitalDelayType01Z := (2 ns,2 ns,2 ns,2 ns,2 ns,2 ns);
tpd_OE_WRDATA0         :VitalDelayType01Z := (2 ns,2 ns,2 ns,2 ns,2 ns,2 ns);
tpd_OE_WRDATA1         :VitalDelayType01Z := (2 ns,2 ns,2 ns,2 ns,2 ns,2 ns);
tpd_OE_WRDATA2         :VitalDelayType01Z := (2 ns,2 ns,2 ns,2 ns,2 ns,2 ns);
tpd_OE_WRDATA3         :VitalDelayType01Z := (2 ns,2 ns,2 ns,2 ns,2 ns,2 ns);
tpd_RAD4_RDATA0         :VitalDelayType01 := (2.0 ns,2.0 ns);
tpd_RAD3_RDATA0         :VitalDelayType01 := (2.0 ns,2.0 ns);
tpd_RAD2_RDATA0         :VitalDelayType01 := (2.0 ns,2.0 ns);
tpd_RAD1_RDATA0         :VitalDelayType01 := (2.0 ns,2.0 ns);
tpd_RAD0_RDATA0         :VitalDelayType01 := (2.0 ns,2.0 ns);
tpd_RAD4_RDATA1         :VitalDelayType01 := (2.0 ns,2.0 ns);
tpd_RAD3_RDATA1         :VitalDelayType01 := (2.0 ns,2.0 ns);
tpd_RAD2_RDATA1         :VitalDelayType01 := (2.0 ns,2.0 ns);
tpd_RAD1_RDATA1         :VitalDelayType01 := (2.0 ns,2.0 ns);
tpd_RAD0_RDATA1         :VitalDelayType01 := (2.0 ns,2.0 ns);
tpd_RAD4_RDATA2         :VitalDelayType01 := (2.0 ns,2.0 ns);
tpd_RAD3_RDATA2         :VitalDelayType01 := (2.0 ns,2.0 ns);
tpd_RAD2_RDATA2         :VitalDelayType01 := (2.0 ns,2.0 ns);
tpd_RAD1_RDATA2         :VitalDelayType01 := (2.0 ns,2.0 ns);
tpd_RAD0_RDATA2         :VitalDelayType01 := (2.0 ns,2.0 ns);
tpd_RAD4_RDATA3         :VitalDelayType01 := (2.0 ns,2.0 ns);
tpd_RAD3_RDATA3         :VitalDelayType01 := (2.0 ns,2.0 ns);
tpd_RAD2_RDATA3         :VitalDelayType01 := (2.0 ns,2.0 ns);
tpd_RAD1_RDATA3         :VitalDelayType01 := (2.0 ns,2.0 ns);
tpd_RAD0_RDATA3         :VitalDelayType01 := (2.0 ns,2.0 ns);

tsetup_WRDATA3_WRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
thold_WRDATA3_WRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
tsetup_WRDATA2_WRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
thold_WRDATA2_WRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
tsetup_WRDATA1_WRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
thold_WRDATA1_WRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
tsetup_WRDATA0_WRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
thold_WRDATA0_WRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
tsetup_WRAD4_WRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
thold_WRAD4_WRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
tsetup_WRAD3_WRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
thold_WRAD3_WRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
tsetup_WRAD2_WRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
thold_WRAD2_WRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
tsetup_WRAD1_WRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
thold_WRAD1_WRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
tsetup_WRAD0_WRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
thold_WRAD0_WRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
tpw_WRCLK_posedge        :VitalDelayType := 1.0 ns;
tsetup_WEN_WRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
thold_WEN_WRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;


        TimingChecksOn : BOOLEAN := TRUE;
	InstancePath : STRING := "*"
            );
  PORT	(
	WEN		: IN	std_logic ;
	REN		: IN	std_logic ;
	WRCLK		: IN	std_logic ;
	OE		: IN	std_logic ;
        WRDATA3         : INOUT std_logic := 'Z';
        WRDATA2         : INOUT std_logic := 'Z';
        WRDATA1         : INOUT std_logic := 'Z';
        WRDATA0         : INOUT std_logic := 'Z';
        RDATA3          :OUT std_logic := 'X';
        RDATA2          : OUT std_logic := 'X';
        RDATA1          : OUT std_logic := 'X';
        RDATA0          : OUT std_logic := 'X';
        RAD4           : IN    std_logic;
        RAD3           : IN    std_logic;
        RAD2           : IN    std_logic;
        RAD1           : IN    std_logic;
        RAD0           : IN    std_logic;
        WRAD4           : IN    std_logic;
        WRAD3           : IN    std_logic;
        WRAD2           : IN    std_logic;
        WRAD1           : IN    std_logic;
        WRAD0           : IN    std_logic
	);


   ATTRIBUTE VITAL_LEVEL0 OF RB_DA : ENTITY IS TRUE;

END RB_DA;

-----------------------------------------------------------------------
-- ARCHITECTURE declaration
-----------------------------------------------------------------------
ARCHITECTURE VITAL_VF OF RB_DA IS

    ATTRIBUTE VITAL_LEVEL1 OF VITAL_VF : ARCHITECTURE IS FALSE;

	SIGNAL WEN_ipd		: std_logic := 'X';
	SIGNAL REN_ipd		: std_logic := 'X';
	SIGNAL WRCLK_ipd		: std_logic := '0';
	SIGNAL WR_CLK		: std_logic := '0';
	SIGNAL OE_ipd	: std_logic := 'X';
        SIGNAL WRDATA3_ipd      : std_logic := 'Z';
        SIGNAL WRDATA2_ipd      : std_logic := 'Z';
        SIGNAL WRDATA1_ipd      : std_logic := 'Z';
        SIGNAL WRDATA0_ipd      : std_logic := 'Z';
        SIGNAL WRAD4_ipd                : std_logic := '0';
        SIGNAL WRAD3_ipd                : std_logic := '0';
        SIGNAL WRAD2_ipd                : std_logic := '0';
        SIGNAL WRAD1_ipd                : std_logic := '0';
        SIGNAL WRAD0_ipd                : std_logic := '0';
        SIGNAL RAD4_ipd                : std_logic := '0';
        SIGNAL RAD3_ipd                : std_logic := '0';
        SIGNAL RAD2_ipd                : std_logic := '0';
        SIGNAL RAD1_ipd                : std_logic := '0';
        SIGNAL RAD0_ipd                : std_logic := '0';
	SIGNAL DIN		: std_logic_vector(3 DOWNTO 0);
	SIGNAL RD_ADD		: std_logic_vector(4 DOWNTO 0);
	SIGNAL RD_ADD_W		: std_logic_vector(4 DOWNTO 0);
	SIGNAL WR_ADD		: std_logic_vector(4 DOWNTO 0);
	SIGNAL write_add	: std_logic_vector(4 DOWNTO 0);
	SIGNAL data_out		: std_logic_vector(3 DOWNTO 0) := x_data;
	SIGNAL data_out_w		: std_logic_vector(3 DOWNTO 0) := z_data;
	SIGNAL output_delay	: time		:= 0 ns;
	SIGNAL output_delay_w	: time		:= 0 ns;
	SIGNAL memory_array	: memory_array_typ;

BEGIN
   
  ---------------------------------------------------------------------
  -- INPUT PATH DELAYs
  ---------------------------------------------------------------------
  WIREDELAY : BLOCK
  BEGIN
	VitalWireDelay (WEN_ipd,		WEN,		tipd_WEN);
	VitalWireDelay (REN_ipd,		REN,		tipd_REN);
	VitalWireDelay (WRCLK_ipd,		WRCLK,		tipd_WRCLK);
	VitalWireDelay (OE_ipd,		OE,		tipd_OE);
        VitalWireDelay (WRDATA0_ipd,    WRDATA0,        tipd_WRDATA0);
        VitalWireDelay (WRDATA1_ipd,    WRDATA1,        tipd_WRDATA1);
        VitalWireDelay (WRDATA2_ipd,    WRDATA2,        tipd_WRDATA2);
        VitalWireDelay (WRDATA3_ipd,    WRDATA3,        tipd_WRDATA3);
        VitalWireDelay (RAD0_ipd,              RAD0,          tipd_RAD0);
        VitalWireDelay (RAD1_ipd,              RAD1,          tipd_RAD1);
        VitalWireDelay (RAD2_ipd,              RAD2,          tipd_RAD2);
        VitalWireDelay (RAD3_ipd,              RAD3,          tipd_RAD3);
        VitalWireDelay (RAD4_ipd,              RAD4,          tipd_RAD4);
        VitalWireDelay (WRAD0_ipd,              WRAD0,          tipd_WRAD0);
        VitalWireDelay (WRAD1_ipd,              WRAD1,          tipd_WRAD1);
        VitalWireDelay (WRAD2_ipd,              WRAD2,          tipd_WRAD2);
        VitalWireDelay (WRAD3_ipd,              WRAD3,          tipd_WRAD3);
        VitalWireDelay (WRAD4_ipd,              WRAD4,          tipd_WRAD4);

  END BLOCK;

  ---------------------------------------------------------------------
  -- Behavior Section
  ---------------------------------------------------------------------

  ---------------------------------------------------------------------
  -- Wrapper Section
  ---------------------------------------------------------------------

   wrapper_read_add : process(REN_ipd, WEN_ipd, OE_ipd, WRAD4_ipd, WRAD3_ipd, WRAD2_ipd, WRAD1_ipd, WRAD0_ipd, RAD4_ipd, RAD3_ipd, RAD2_ipd, RAD1_ipd, RAD0_ipd)

   begin
    if (REN_ipd = '1') then
        RD_ADD(4) <= RAD4_ipd;
        RD_ADD(3) <= RAD3_ipd;
        RD_ADD(2) <= RAD2_ipd;
        RD_ADD(1) <= RAD1_ipd;
        RD_ADD(0) <= RAD0_ipd;
    else
	RD_ADD <= x_add;
    end if;

    if (REN_ipd = '1' and WEN_ipd = '0' and OE_ipd = '1') then
        RD_ADD_W(4) <= WRAD4_ipd;
        RD_ADD_W(3) <= WRAD3_ipd;
        RD_ADD_W(2) <= WRAD2_ipd;
        RD_ADD_W(1) <= WRAD1_ipd;
        RD_ADD_W(0) <= WRAD0_ipd;
    else
	RD_ADD_W <= x_add;
    end if;

   end process;

   wrapper_write_add : process(WEN_ipd, WRAD4_ipd, WRAD3_ipd, WRAD2_ipd, WRAD1_ipd, WRAD0_ipd)

   begin
    if (WEN_ipd = '1') then
        WR_ADD(4) <= WRAD4_ipd;
        WR_ADD(3) <= WRAD3_ipd;
        WR_ADD(2) <= WRAD2_ipd;
        WR_ADD(1) <= WRAD1_ipd;
        WR_ADD(0) <= WRAD0_ipd;
    else
	WR_ADD <= x_add;
    end if;

   end process;

   wrapper_write_clk : process(WEN_ipd, WRCLK_ipd)

   begin
    if (WEN_ipd = '1') then
	WR_CLK <= WRCLK_ipd;
    else
	WR_CLK <= '0';
    end if;

   end process;

   process(WR_CLK)

    begin
      if WR_CLK = '1' then
        write_add(4) <= WRAD4_ipd;
        write_add(3) <= WRAD3_ipd;
        write_add(2) <= WRAD2_ipd;
        write_add(1) <= WRAD1_ipd;
        write_add(0) <= WRAD0_ipd;
      end if;

   end process;

   wrapper_write_data : process(WEN_ipd, WRDATA3_ipd, WRDATA2_ipd, WRDATA1_ipd, WRDATA0_ipd)

   begin
    if (WEN_ipd = '1') then
        DIN(3) <= WRDATA3_ipd;
        DIN(2) <= WRDATA2_ipd;
        DIN(1) <= WRDATA1_ipd;
        DIN(0) <= WRDATA0_ipd;
    else
	DIN <= x_data;
    end if;

   end process;


  VITALBehavior : PROCESS ( WEN_ipd, REN_ipd, WR_CLK,  DIN, RD_ADD_W, RD_ADD, WR_ADD,  RAD4_ipd, RAD3_ipd, RAD2_ipd, RAD1_ipd, RAD0_ipd, WRAD4_ipd,WRAD3_ipd,WRAD2_ipd,WRAD1_ipd,WRAD0_ipd )


   -- Temporary variables
   VARIABLE tempaddr 		: integer := 0;
   VARIABLE rd_address 		: integer := 0;
   VARIABLE rd_address_w 	: integer := 0;

   -- Timing Check results
   VARIABLE Pviol_WRCLK			: std_logic := '0';
   VARIABLE PeriodData_WRCLK		: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_WR_ADD_stp_hld_0	: std_logic := '0';
   VARIABLE TimingData_WR_ADD_stp_hld_0	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_WR_ADD_stp_hld_1	: std_logic := '0';
   VARIABLE TimingData_WR_ADD_stp_hld_1	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_WR_ADD_stp_hld_2	: std_logic := '0';
   VARIABLE TimingData_WR_ADD_stp_hld_2	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_WR_ADD_stp_hld_3	: std_logic := '0';
   VARIABLE TimingData_WR_ADD_stp_hld_3	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_WR_ADD_stp_hld_4	: std_logic := '0';
   VARIABLE TimingData_WR_ADD_stp_hld_4	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_WR_DATA_stp_0		: std_logic := '0';
   VARIABLE TimingData_WR_DATA_stp_0	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_WR_DATA_stp_1		: std_logic := '0';
   VARIABLE TimingData_WR_DATA_stp_1	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_WR_DATA_stp_2		: std_logic := '0';
   VARIABLE TimingData_WR_DATA_stp_2	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_WR_DATA_stp_3		: std_logic := '0';
   VARIABLE TimingData_WR_DATA_stp_3	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_WR_DATA_hld_0		: std_logic := '0';
   VARIABLE TimingData_WR_DATA_hld_0	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_WR_DATA_hld_1		: std_logic := '0';
   VARIABLE TimingData_WR_DATA_hld_1	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_WR_DATA_hld_2		: std_logic := '0';
   VARIABLE TimingData_WR_DATA_hld_2	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_WR_DATA_hld_3		: std_logic := '0';
   VARIABLE TimingData_WR_DATA_hld_3	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_WEN_hld		: std_logic := '0';
   VARIABLE TimingData_WEN_hld		: VitalTimingDataType := VitalTimingDataInit;



 BEGIN
    -------------------------------------------------------------------
    -- Timing Check Section
    -------------------------------------------------------------------
    IF (TimingChecksOn) THEN

        VitalPeriodPulseCheck  (Pviol_WRCLK,
                                PeriodData_WRCLK,
                                WR_CLK, "WRCLK",
                                0.0 ns,
                                0.0 ns,
                                tpw_WRCLK_posedge,
                                0.0 ns,
                                TRUE,
                                InstancePath & "/RB_DA",
                                TRUE,
                                TRUE,
                                WARNING );

        VitalSetupHoldCheck    (Tviol_WR_ADD_stp_hld_0,
                                TimingData_WR_ADD_stp_hld_0,
                                WR_ADD(0), "WRAD0",
                                0.0 ns,
                                WR_CLK, "WRCLK",
                                0.0 ns,
                                tsetup_WRAD0_WRCLK_noedge_posedge, tsetup_WRAD0_WRCLK_noedge_posedge,
                                thold_WRAD0_WRCLK_noedge_posedge, thold_WRAD0_WRCLK_noedge_posedge,
                                WEN_ipd = '1',
                                '/',
                                InstancePath & "/RB_DA",
                                TRUE,
                                TRUE,
                                WARNING );

        VitalSetupHoldCheck    (Tviol_WR_ADD_stp_hld_1,
                                TimingData_WR_ADD_stp_hld_1,
                                WR_ADD(1), "WRAD1",
                                0.0 ns,
                                WR_CLK, "WRCLK",
                                0.0 ns,
                                tsetup_WRAD1_WRCLK_noedge_posedge, tsetup_WRAD1_WRCLK_noedge_posedge,
                                thold_WRAD1_WRCLK_noedge_posedge, thold_WRAD1_WRCLK_noedge_posedge,
                                WEN_ipd = '1',
                                '/',
                                InstancePath & "/RB_DA",
                                TRUE,
                                TRUE,
                                WARNING );

        VitalSetupHoldCheck    (Tviol_WR_ADD_stp_hld_2,
                                TimingData_WR_ADD_stp_hld_2,
                                WR_ADD(2), "WRAD2",
                                0.0 ns,
                                WR_CLK, "WRCLK",
                                0.0 ns,
                                tsetup_WRAD2_WRCLK_noedge_posedge, tsetup_WRAD2_WRCLK_noedge_posedge,
                                thold_WRAD2_WRCLK_noedge_posedge, thold_WRAD2_WRCLK_noedge_posedge,
                                WEN_ipd = '1',
                                '/',
                                InstancePath & "/RB_DA",
                                TRUE,
                                TRUE,
                                WARNING );
       VitalSetupHoldCheck    (Tviol_WR_ADD_stp_hld_3,
                                TimingData_WR_ADD_stp_hld_3,
                                WR_ADD(3), "WRAD3",
                                0.0 ns,
                                WR_CLK, "WRCLK",
                                0.0 ns,
                                tsetup_WRAD3_WRCLK_noedge_posedge, tsetup_WRAD3_WRCLK_noedge_posedge,
                                thold_WRAD3_WRCLK_noedge_posedge, thold_WRAD3_WRCLK_noedge_posedge,
                                WEN_ipd = '1',
                                '/',
                                InstancePath & "/RB_DA",
                                TRUE,
                                TRUE,
                                WARNING );
        VitalSetupHoldCheck    (Tviol_WR_ADD_stp_hld_4,
                                TimingData_WR_ADD_stp_hld_4,
                                WR_ADD(4), "WRAD4",
                                0.0 ns,
                                WR_CLK, "WRCLK",
                                0.0 ns,
                                tsetup_WRAD4_WRCLK_noedge_posedge, tsetup_WRAD4_WRCLK_noedge_posedge,
                                thold_WRAD4_WRCLK_noedge_posedge, thold_WRAD4_WRCLK_noedge_posedge,
                                WEN_ipd = '1',
                                '/',
                                InstancePath & "/RB_DA",
                                TRUE,
                                TRUE,
                                WARNING );

        VitalSetupHoldCheck    (Tviol_WR_DATA_stp_0,
                                TimingData_WR_DATA_stp_0,
                                DIN(0), "WRDATA0",
                                0.0 ns,
                                WR_CLK, "WRCLK",
                                0.0 ns,
                                tsetup_WRDATA0_WRCLK_noedge_posedge, tsetup_WRDATA0_WRCLK_noedge_posedge,
                                0.0 ns, 0.0 ns,
                                WEN_ipd = '1',
                                '/',
                                InstancePath & "/RB_DA",
                                TRUE,
                                TRUE,
                                WARNING );

        VitalSetupHoldCheck    (Tviol_WR_DATA_stp_1,
                                TimingData_WR_DATA_stp_1,
                                DIN(1), "WRDATA1",
                                0.0 ns,
                                WR_CLK, "WRCLK",
                                0.0 ns,
                                tsetup_WRDATA1_WRCLK_noedge_posedge, tsetup_WRDATA1_WRCLK_noedge_posedge,
                                0.0 ns, 0.0 ns,
                                WEN_ipd = '1',
                                '/',
                                InstancePath & "/RB_DA",
                                TRUE,
                                TRUE,
                                WARNING );

        VitalSetupHoldCheck    (Tviol_WR_DATA_stp_2,
                                TimingData_WR_DATA_stp_2,
                                DIN(2), "WRDATA2",
                                0.0 ns,
                                WR_CLK, "WRCLK",
                                0.0 ns,
                                tsetup_WRDATA2_WRCLK_noedge_posedge, tsetup_WRDATA2_WRCLK_noedge_posedge,
                                0.0 ns, 0.0 ns,
                                WEN_ipd = '1',
                                '/',
                                InstancePath & "/RB_DA",
                                TRUE,
                                TRUE,
                                WARNING );

        VitalSetupHoldCheck    (Tviol_WR_DATA_stp_3,
                                TimingData_WR_DATA_stp_3,
                                DIN(3), "WRDATA3",
                                0.0 ns,
                                WR_CLK, "WRCLK",
                                0.0 ns,
                                tsetup_WRDATA3_WRCLK_noedge_posedge, tsetup_WRDATA3_WRCLK_noedge_posedge,
                                0.0 ns, 0.0 ns,
                                WEN_ipd = '1',
                                '/',
                                InstancePath & "/RB_DA",
                                TRUE,
                                TRUE,
                                WARNING );

        VitalSetupHoldCheck    (Tviol_WR_DATA_hld_0,
                                TimingData_WR_DATA_hld_0,
                                DIN(0), "WRDATA0",
                                0.0 ns,
                                WR_CLK, "WRCLK",
                                0.0 ns,
                                0.0 ns, 0.0 ns,
                                thold_WRDATA0_WRCLK_noedge_posedge, thold_WRDATA0_WRCLK_noedge_posedge,
                                WEN_ipd = '1',
                                '/',
                                InstancePath & "/RB_DA",
                                TRUE,
                                TRUE,
                                WARNING );

        VitalSetupHoldCheck    (Tviol_WR_DATA_hld_1,
                                TimingData_WR_DATA_hld_1,
                                DIN(1), "WRDATA1",
                                0.0 ns,
                                WR_CLK, "WRCLK",
                                0.0 ns,
                                0.0 ns, 0.0 ns,
                                thold_WRDATA1_WRCLK_noedge_posedge, thold_WRDATA1_WRCLK_noedge_posedge,
                                WEN_ipd = '1',
                                '/',
                                InstancePath & "/RB_DA",
                                TRUE,
                                TRUE,
                                WARNING );

        VitalSetupHoldCheck    (Tviol_WR_DATA_hld_2,
                                TimingData_WR_DATA_hld_2,
                                DIN(2), "WRDATA2",
                                0.0 ns,
                                WR_CLK, "WRCLK",
                                0.0 ns,
                                0.0 ns, 0.0 ns,
                                thold_WRDATA2_WRCLK_noedge_posedge, thold_WRDATA2_WRCLK_noedge_posedge,
                                WEN_ipd = '1',
                                '/',
                                InstancePath & "/RB_DA",
                                TRUE,
                                TRUE,
                                WARNING );
        VitalSetupHoldCheck    (Tviol_WR_DATA_hld_3,
                                TimingData_WR_DATA_hld_3,
                                DIN(3), "WRDATA3",
                                0.0 ns,
                                WR_CLK, "WRCLK",
                                0.0 ns,
                                0.0 ns, 0.0 ns,
                                thold_WRDATA3_WRCLK_noedge_posedge, thold_WRDATA3_WRCLK_noedge_posedge,
                                WEN_ipd = '1',
                                '/',
                                InstancePath & "/RB_DA",
                                TRUE,
                                TRUE,
                                WARNING );


        VitalSetupHoldCheck    (Tviol_WEN_hld,
                                TimingData_WEN_hld,
                                WEN_ipd, "WEN",
                                0.0 ns,
                                WR_CLK, "WRCLK",
                                0.0 ns,
                                tsetup_WEN_WRCLK_noedge_posedge, tsetup_WEN_WRCLK_noedge_posedge,
                                thold_WEN_WRCLK_noedge_posedge, thold_WEN_WRCLK_noedge_posedge,
                                True,
                                '/',
                                InstancePath & "/RB_DA",
                                TRUE,
                                TRUE,
                                WARNING );

    END IF; -- Timing Check Section

    -------------------------------------------------------------------
    -- Functionality Section
    -------------------------------------------------------------------

-- WRITE ADDRESS GOES XX

    if ( WR_CLK'EVENT and WR_CLK = '1' and vecX(WR_ADD)) then

        assert false
        report "Illegal Address Input: Undefined  Address at the Read_Write Port."
        severity note ;
        memory_array <= (others => x_data);

    end if;

-- ADDRESS HOLD AND SETUP VIOLATION EFFECT

    if( Tviol_WR_ADD_stp_hld_0 = 'X' or Tviol_WR_ADD_stp_hld_1 = 'X' or Tviol_WR_ADD_stp_hld_2 = 'X' or Tviol_WR_ADD_stp_hld_3 = 'X' or Tviol_WR_ADD_stp_hld_4 = 'X' ) then

        memory_array <= (others => x_data);

    else

-- DATA SETUP AND HOLD VIOLATION EFFECT

    if( Pviol_WRCLK = 'X' or Tviol_WR_DATA_hld_0 = 'X' or Tviol_WR_DATA_hld_1 = 'X' or Tviol_WR_DATA_hld_2 = 'X' or Tviol_WR_DATA_hld_3 = 'X' or Tviol_WEN_hld = 'X') then
	tempaddr := vec2int(write_add);
	memory_array(tempaddr) <= x_data;
    end if;

    if( Tviol_WR_DATA_stp_0 = 'X' or Tviol_WR_DATA_stp_1 = 'X' or Tviol_WR_DATA_stp_2 = 'X' or Tviol_WR_DATA_stp_3 = 'X') then
	tempaddr := vec2int(WR_ADD);
	memory_array(tempaddr) <= x_data;
    end if;

    end if;

-- VALID MEMORY WRITE

    if ( WR_CLK'EVENT and WR_CLK = '1' and not(vecX(WR_ADD)) and not(Tviol_WR_ADD_stp_hld_0 = 'X' or Tviol_WR_ADD_stp_hld_1 = 'X' or Tviol_WR_ADD_stp_hld_2 = 'X' or Tviol_WR_ADD_stp_hld_3 = 'X' or Tviol_WR_ADD_stp_hld_4 = 'X') and not( Pviol_WRCLK = 'X' or Tviol_WR_DATA_hld_0 = 'X' or Tviol_WR_DATA_hld_1 = 'X' or Tviol_WR_DATA_hld_2 = 'X' or Tviol_WR_DATA_hld_3 = 'X' or Tviol_WEN_hld = 'X') and not( Tviol_WR_DATA_stp_0 = 'X' or Tviol_WR_DATA_stp_1 = 'X' or Tviol_WR_DATA_stp_2 = 'X' or Tviol_WR_DATA_stp_3 = 'X')) then
	tempaddr := vec2int(WR_ADD);
	memory_array(tempaddr) <= DIN;
    end if;

    if WR_CLK'EVENT and WR_CLK /= WRCLK_ipd and WR_CLK'LAST_VALUE = '1' then
	memory_array(tempaddr) <= x_data;
    end if;


-- READ CYCLE VIOLATION EFFECT

    if(RD_ADD'EVENT and REN_ipd = '1' and vecX(RD_ADD)) then
	data_out <= x_data;
    elsif

-- VALID MEMORY READ

     (RD_ADD'EVENT and REN_ipd = '1'  and not (vecX(RD_ADD))) then
	rd_address := vec2int(RD_ADD);
	data_out <= memory_array(rd_address);
    end if;

    if(RD_ADD_W'EVENT and REN_ipd = '1' and OE_ipd = '1' and vecX(RD_ADD_W)) then
	data_out_w <= x_data;
    elsif

-- VALID MEMORY READ

     (RD_ADD_W'EVENT  and REN_ipd = '1' and OE_ipd = '1' and WEN_ipd = '0' and not (vecX(RD_ADD_W))) then
	rd_address_w := vec2int(RD_ADD_W);
	data_out_w <= memory_array(rd_address_w);
    end if;

  END PROCESS;

    -------------------------------------------------------------------------------
    -- Temporary output signal should get assigned to the output signal.
    -------------------------------------------------------------------------------

   PROCESS(data_out, data_out_w, REN_ipd, OE_ipd, RAD4_ipd, RAD3_ipd, RAD2_ipd, RAD1_ipd, RAD0_ipd, WRAD4_ipd, WRAD3_ipd, WRAD2_ipd, WRAD1_ipd, WRAD0_ipd)

   VARIABLE GLITCH_DATA : VitalGlitchDataType;
   VARIABLE GLITCH : VitalGlitchDataType;
   VARIABLE con : std_logic ;--:= '0';
    VARIABLE WEN_inv : std_logic ;--:= '0';
    VARIABLE WRDATA3_1 : std_logic := 'Z';
    VARIABLE WRDATA2_1 : std_logic := 'Z';
    VARIABLE WRDATA1_1 : std_logic := 'Z';
    VARIABLE WRDATA0_1 : std_logic := 'Z';
    VARIABLE RDATA3_1 : std_logic := 'X';
    VARIABLE RDATA2_1 : std_logic := 'X';
    VARIABLE RDATA1_1 : std_logic := 'X';
    VARIABLE RDATA0_1 : std_logic := 'X';

   BEGIN
       WEN_inv := VitalINV(WEN_ipd);
       con := VitalAND3(OE_ipd,REN_ipd, WEN_inv);


      WRDATA3_1 := VITALBUFIF1(data_out_w(3),con);
      WRDATA2_1 := VITALBUFIF1(data_out_w(2),con);
      WRDATA1_1 := VITALBUFIF1(data_out_w(1),con);
      WRDATA0_1 := VITALBUFIF1(data_out_w(0),con);

      RDATA3_1 := VITALBUF(data_out(3));
      RDATA2_1 := VITALBUF(data_out(2));
      RDATA1_1 := VITALBUF(data_out(1));
      RDATA0_1 := VITALBUF(data_out(0));

     VitalPathDelay01 ( RDATA3, GLITCH, "RDATA3", RDATA3_1,
        Paths => (
        0 => ( RAD4_ipd'LAST_EVENT, tpd_RAD4_RDATA3, TRUE ),
        1 => ( RAD3_ipd'LAST_EVENT, tpd_RAD3_RDATA3, TRUE ),
        2 => ( RAD2_ipd'LAST_EVENT, tpd_RAD2_RDATA3, TRUE ),
        3 => ( RAD1_ipd'LAST_EVENT, tpd_RAD1_RDATA3, TRUE ),
        4 => ( RAD0_ipd'LAST_EVENT, tpd_RAD0_RDATA3, TRUE )),
        DefaultDelay=>VitalZeroDelay01,
        Mode=>VitalInertial,
        XON=>TRUE,
        MsgOn=>TRUE,
        MsgSeverity=>WARNING );

     VitalPathDelay01 ( RDATA2, GLITCH, "RDATA2", RDATA2_1,
        Paths => (
        0 => ( RAD4_ipd'LAST_EVENT, tpd_RAD4_RDATA2, TRUE ),
        1 => ( RAD3_ipd'LAST_EVENT, tpd_RAD3_RDATA2, TRUE ),
        2 => ( RAD2_ipd'LAST_EVENT, tpd_RAD2_RDATA2, TRUE ),
        3 => ( RAD1_ipd'LAST_EVENT, tpd_RAD1_RDATA2, TRUE ),
        4 => ( RAD0_ipd'LAST_EVENT, tpd_RAD0_RDATA2, TRUE )),
        DefaultDelay=>VitalZeroDelay01,
        Mode=>VitalInertial,
        XON=>TRUE,
        MsgOn=>TRUE,
        MsgSeverity=>WARNING );

     VitalPathDelay01 ( RDATA1, GLITCH, "RDATA1", RDATA1_1,
        Paths => (
        0 => ( RAD4_ipd'LAST_EVENT, tpd_RAD4_RDATA1, TRUE ),
        1 => ( RAD3_ipd'LAST_EVENT, tpd_RAD3_RDATA1, TRUE ),
        2 => ( RAD2_ipd'LAST_EVENT, tpd_RAD2_RDATA1, TRUE ),
        3 => ( RAD1_ipd'LAST_EVENT, tpd_RAD1_RDATA1, TRUE ),
        4 => ( RAD0_ipd'LAST_EVENT, tpd_RAD0_RDATA1, TRUE )),
        DefaultDelay=>VitalZeroDelay01,
        Mode=>VitalInertial,
        XON=>TRUE,
        MsgOn=>TRUE,
        MsgSeverity=>WARNING );

     VitalPathDelay01 ( RDATA0, GLITCH, "RDATA0", RDATA0_1,
        Paths => (
        0 => ( RAD4_ipd'LAST_EVENT, tpd_RAD4_RDATA0, TRUE ),
        1 => ( RAD3_ipd'LAST_EVENT, tpd_RAD3_RDATA0, TRUE ),
        2 => ( RAD2_ipd'LAST_EVENT, tpd_RAD2_RDATA0, TRUE ),
        3 => ( RAD1_ipd'LAST_EVENT, tpd_RAD1_RDATA0, TRUE ),
        4 => ( RAD0_ipd'LAST_EVENT, tpd_RAD0_RDATA0, TRUE )),
        DefaultDelay=>VitalZeroDelay01,
        Mode=>VitalInertial,
        XON=>TRUE,
        MsgOn=>TRUE,
        MsgSeverity=>WARNING );


      VitalPathDelay01Z ( WRDATA3, GLITCH_DATA, "WRDATA3", WRDATA3_1,
        Paths => (
        0 => ( WRAD4_ipd'LAST_EVENT, VitalExtendToFillDelay(tpd_WRAD4_WRDATA3), TRUE ),
        1 => ( WRAD3_ipd'LAST_EVENT, VitalExtendToFillDelay(tpd_WRAD3_WRDATA3), TRUE ),
        2 => ( WRAD2_ipd'LAST_EVENT, VitalExtendToFillDelay(tpd_WRAD2_WRDATA3), TRUE ),
        3 => ( WRAD1_ipd'LAST_EVENT, VitalExtendToFillDelay(tpd_WRAD1_WRDATA3), TRUE ),
        4 => ( WRAD0_ipd'LAST_EVENT, VitalExtendToFillDelay(tpd_WRAD0_WRDATA3), TRUE ),
        5 => ( OE_ipd'LAST_EVENT, VitalExtendToFillDelay(tpd_OE_WRDATA3), TRUE ) ),
        DefaultDelay=>VitalZeroDelay01Z,
        Mode=>VitalInertial,
        XON=>TRUE,
        MsgOn=>TRUE,
        MsgSeverity=>WARNING,
        OutputMap => "UX01ZWLH-");

      VitalPathDelay01Z ( WRDATA2, GLITCH_DATA, "WRDATA2", WRDATA2_1,
        Paths => (
        0 => ( WRAD4_ipd'LAST_EVENT, VitalExtendToFillDelay(tpd_WRAD4_WRDATA2), TRUE ),
        1 => ( WRAD3_ipd'LAST_EVENT, VitalExtendToFillDelay(tpd_WRAD3_WRDATA2), TRUE ),
        2 => ( WRAD2_ipd'LAST_EVENT, VitalExtendToFillDelay(tpd_WRAD2_WRDATA2), TRUE ),
        3 => ( WRAD1_ipd'LAST_EVENT, VitalExtendToFillDelay(tpd_WRAD1_WRDATA2), TRUE ),
        4 => ( WRAD0_ipd'LAST_EVENT, VitalExtendToFillDelay(tpd_WRAD0_WRDATA2), TRUE ),
        5 => ( OE_ipd'LAST_EVENT, VitalExtendToFillDelay(tpd_OE_WRDATA2), TRUE ) ),
        DefaultDelay=>VitalZeroDelay01Z,
        Mode=>VitalInertial,
        XON=>TRUE,
        MsgOn=>TRUE,
        MsgSeverity=>WARNING,
        OutputMap => "UX01ZWLH-");

      VitalPathDelay01Z ( WRDATA1, GLITCH_DATA, "WRDATA1", WRDATA1_1,
        Paths => (
        0 => ( WRAD4_ipd'LAST_EVENT, VitalExtendToFillDelay(tpd_WRAD4_WRDATA1), TRUE ),
        1 => ( WRAD3_ipd'LAST_EVENT, VitalExtendToFillDelay(tpd_WRAD3_WRDATA1), TRUE ),
        2 => ( WRAD2_ipd'LAST_EVENT, VitalExtendToFillDelay(tpd_WRAD2_WRDATA1), TRUE ),
        3 => ( WRAD1_ipd'LAST_EVENT, VitalExtendToFillDelay(tpd_WRAD1_WRDATA1), TRUE ),
        4 => ( WRAD0_ipd'LAST_EVENT, VitalExtendToFillDelay(tpd_WRAD0_WRDATA1), TRUE ),
        5 => ( OE_ipd'LAST_EVENT, VitalExtendToFillDelay(tpd_OE_WRDATA1), TRUE ) ),
        DefaultDelay=>VitalZeroDelay01Z,
        Mode=>VitalInertial,
        XON=>TRUE,
        MsgOn=>TRUE,
        MsgSeverity=>WARNING,
        OutputMap => "UX01ZWLH-");

       VitalPathDelay01Z ( WRDATA0, GLITCH_DATA, "WRDATA0", WRDATA0_1,
        Paths => (
        0 => ( WRAD4_ipd'LAST_EVENT, VitalExtendToFillDelay(tpd_WRAD4_WRDATA0), TRUE ),
        1 => ( WRAD3_ipd'LAST_EVENT, VitalExtendToFillDelay(tpd_WRAD3_WRDATA0), TRUE ),
        2 => ( WRAD2_ipd'LAST_EVENT, VitalExtendToFillDelay(tpd_WRAD2_WRDATA0), TRUE ),
        3 => ( WRAD1_ipd'LAST_EVENT, VitalExtendToFillDelay(tpd_WRAD1_WRDATA0), TRUE ),
        4 => ( WRAD0_ipd'LAST_EVENT, VitalExtendToFillDelay(tpd_WRAD0_WRDATA0), TRUE ),
        5 => ( OE_ipd'LAST_EVENT, VitalExtendToFillDelay(tpd_OE_WRDATA0), TRUE ) ),
        DefaultDelay=>VitalZeroDelay01Z,
        Mode=>VitalInertial,
        XON=>TRUE,
        MsgOn=>TRUE,
        MsgSeverity=>WARNING,
        OutputMap => "UX01ZWLH-");

END PROCESS;



END VITAL_VF;
configuration CFG_RB_DA_VITAL of RB_DA is
        for VITAL_VF
        end for;
end CFG_RB_DA_VITAL;
-----------------------------------------------------------------------


-----------------------------------------------------------------------
-- VITAL model for RB_DS 30.10 technology
-----------------------------------------------------------------------

LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.VITAL_timing.all;
USE IEEE.VITAL_primitives.all;
LIBRARY VF1;
USE VF1.ALL;
USE VF1.RAMPACK.ALL;

-----------------------------------------------------------------------
-- ENTITY declaration
-----------------------------------------------------------------------

ENTITY RB_DS IS
  GENERIC (
	tipd_WEN		: VitalDelayType01			:= (0.0 ns, 0.0 ns);
	tipd_REN		: VitalDelayType01			:= (0.0 ns, 0.0 ns);
	tipd_WRCLK		: VitalDelayType01			:= (0.0 ns, 0.0 ns);
	tipd_RCLK		: VitalDelayType01			:= (0.0 ns, 0.0 ns);
	tipd_OE		: VitalDelayType01			:= (0.0 ns, 0.0 ns);
        tipd_WRDATA3            : VitalDelayType01      := (0.0 ns, 0.0 ns);
        tipd_WRDATA2            : VitalDelayType01      := (0.0 ns, 0.0 ns);
        tipd_WRDATA1            : VitalDelayType01      := (0.0 ns, 0.0 ns);
        tipd_WRDATA0            : VitalDelayType01      := (0.0 ns, 0.0 ns);
        tipd_WRAD4              : VitalDelayType01      := (0.0 ns, 0.0 ns);
        tipd_WRAD3              : VitalDelayType01      := (0.0 ns, 0.0 ns);
        tipd_WRAD2              : VitalDelayType01      := (0.0 ns, 0.0 ns);
        tipd_WRAD1              : VitalDelayType01      := (0.0 ns, 0.0 ns);
        tipd_WRAD0              : VitalDelayType01      := (0.0 ns, 0.0 ns);
        tipd_RAD4              : VitalDelayType01      := (0.0 ns, 0.0 ns);
        tipd_RAD3              : VitalDelayType01      := (0.0 ns, 0.0 ns);
        tipd_RAD2              : VitalDelayType01      := (0.0 ns, 0.0 ns);
        tipd_RAD1              : VitalDelayType01      := (0.0 ns, 0.0 ns);
        tipd_RAD0              : VitalDelayType01      := (0.0 ns, 0.0 ns);

tpd_RCLK_RDATA0         :VitalDelayType01 := (2.0 ns,2.0 ns);
tpd_RCLK_RDATA1         :VitalDelayType01 := (2.0 ns,2.0 ns);
tpd_RCLK_RDATA2         :VitalDelayType01 := (2.0 ns,2.0 ns);
tpd_RCLK_RDATA3         :VitalDelayType01 := (2.0 ns,2.0 ns);
tpd_WRCLK_WRDATA0         :VitalDelayType01Z := (2 ns,2 ns,2 ns,2 ns,2 ns,2 ns);
tpd_WRCLK_WRDATA1         :VitalDelayType01Z := (2 ns,2 ns,2 ns,2 ns,2 ns,2 ns);
tpd_WRCLK_WRDATA2         :VitalDelayType01Z := (2 ns,2 ns,2 ns,2 ns,2 ns,2 ns);
tpd_WRCLK_WRDATA3         :VitalDelayType01Z := (2 ns,2 ns,2 ns,2 ns,2 ns,2 ns);
tpd_OE_WRDATA0         :VitalDelayType01Z := (2 ns,2 ns,2 ns,2 ns,2 ns,2 ns);
tpd_OE_WRDATA1         :VitalDelayType01Z := (2 ns,2 ns,2 ns,2 ns,2 ns,2 ns);
tpd_OE_WRDATA2         :VitalDelayType01Z := (2 ns,2 ns,2 ns,2 ns,2 ns,2 ns);
tpd_OE_WRDATA3         :VitalDelayType01Z := (2 ns,2 ns,2 ns,2 ns,2 ns,2 ns);
tpw_WRCLK_posedge        :VitalDelayType := 1.0 ns;
tpw_RCLK_posedge        :VitalDelayType := 1.0 ns;
tsetup_WRDATA3_WRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
thold_WRDATA3_WRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
tsetup_WRDATA2_WRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
thold_WRDATA2_WRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
tsetup_WRDATA1_WRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
thold_WRDATA1_WRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
tsetup_WRDATA0_WRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
thold_WRDATA0_WRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
tsetup_WRAD4_WRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
thold_WRAD4_WRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
tsetup_WRAD3_WRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
thold_WRAD3_WRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
tsetup_WRAD2_WRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
thold_WRAD2_WRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
tsetup_WRAD1_WRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
thold_WRAD1_WRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
tsetup_WRAD0_WRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
thold_WRAD0_WRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
tsetup_WEN_WRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
thold_WEN_WRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
tsetup_RAD4_RCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
thold_RAD4_RCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
tsetup_RAD3_RCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
thold_RAD3_RCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
tsetup_RAD2_RCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
thold_RAD2_RCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
tsetup_RAD1_RCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
thold_RAD1_RCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
tsetup_RAD0_RCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
thold_RAD0_RCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
tsetup_REN_RCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
thold_REN_RCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
	TimingChecksOn : BOOLEAN := TRUE;
	InstancePath : STRING := "*"
            );
  PORT	(
	WEN		: IN	std_logic ;
	REN		: IN	std_logic ;
	WRCLK		: IN	std_logic ;
	RCLK		: IN	std_logic ;
	OE		: IN	std_logic ;
        WRDATA3         : INOUT std_logic := 'Z';
        WRDATA2         : INOUT std_logic := 'Z';
        WRDATA1         : INOUT std_logic := 'Z';
        WRDATA0         : INOUT std_logic := 'Z';
        RDATA3          :OUT std_logic := 'X';
        RDATA2          : OUT std_logic := 'X';
        RDATA1          : OUT std_logic := 'X';
        RDATA0          : OUT std_logic := 'X';
        RAD4           : IN    std_logic;
        RAD3           : IN    std_logic;
        RAD2           : IN    std_logic;
        RAD1           : IN    std_logic;
        RAD0           : IN    std_logic;
        WRAD4           : IN    std_logic;
        WRAD3           : IN    std_logic;
        WRAD2           : IN    std_logic;
        WRAD1           : IN    std_logic;
        WRAD0           : IN    std_logic
	);


   ATTRIBUTE VITAL_LEVEL0 OF RB_DS : ENTITY IS TRUE;

END RB_DS;

-----------------------------------------------------------------------
-- ARCHITECTURE declaration
-----------------------------------------------------------------------
ARCHITECTURE VITAL_VF OF RB_DS IS

    ATTRIBUTE VITAL_LEVEL1 OF VITAL_VF : ARCHITECTURE IS FALSE;

	SIGNAL WEN_ipd		: std_logic := 'X';
	SIGNAL REN_ipd		: std_logic := 'X';
	SIGNAL WRCLK_ipd		: std_logic := '0';
	SIGNAL WR_CLK		: std_logic := '0';
	SIGNAL RCLK_ipd		: std_logic := '0';
	SIGNAL RD_CLK		: std_logic := '0';
	SIGNAL RD_CLK_W		: std_logic := '0';
	SIGNAL OE_ipd	: std_logic := 'X';
	SIGNAL DIN		: std_logic_vector(3 DOWNTO 0);
	SIGNAL RD_ADD		: std_logic_vector(4 DOWNTO 0);
	SIGNAL RD_ADD_W		: std_logic_vector(4 DOWNTO 0);
	SIGNAL WR_ADD		: std_logic_vector(4 DOWNTO 0);
        SIGNAL WRDATA3_ipd      : std_logic := 'Z';
        SIGNAL WRDATA2_ipd      : std_logic := 'Z';
        SIGNAL WRDATA1_ipd      : std_logic := 'Z';
        SIGNAL WRDATA0_ipd      : std_logic := 'Z';
        SIGNAL WRAD4_ipd                : std_logic := '0';
        SIGNAL WRAD3_ipd                : std_logic := '0';
        SIGNAL WRAD2_ipd                : std_logic := '0';
        SIGNAL WRAD1_ipd                : std_logic := '0';
        SIGNAL WRAD0_ipd                : std_logic := '0';
        SIGNAL RAD4_ipd                : std_logic := '0';
        SIGNAL RAD3_ipd                : std_logic := '0';
        SIGNAL RAD2_ipd                : std_logic := '0';
        SIGNAL RAD1_ipd                : std_logic := '0';
        SIGNAL RAD0_ipd                : std_logic := '0';
	SIGNAL write_add	: std_logic_vector(4 DOWNTO 0);
	SIGNAL data_out		: std_logic_vector(3 DOWNTO 0) := x_data;
	SIGNAL data_out_w	: std_logic_vector(3 DOWNTO 0) := z_data;
	SIGNAL output_delay_w	: time		:= 0 ns;
	SIGNAL output_delay	: time		:= 0 ns;

BEGIN
   
  ---------------------------------------------------------------------
  -- INPUT PATH DELAYs
  ---------------------------------------------------------------------
  WIREDELAY : BLOCK
  BEGIN
	VitalWireDelay (WEN_ipd,		WEN,		tipd_WEN);
	VitalWireDelay (REN_ipd,		REN,		tipd_REN);
	VitalWireDelay (WRCLK_ipd,		WRCLK,		tipd_WRCLK);
	VitalWireDelay (RCLK_ipd,		RCLK,		tipd_RCLK);
	VitalWireDelay (OE_ipd,		OE,		tipd_OE);
        VitalWireDelay (WRDATA0_ipd,    WRDATA0,        tipd_WRDATA0);
        VitalWireDelay (WRDATA1_ipd,    WRDATA1,        tipd_WRDATA1);
        VitalWireDelay (WRDATA2_ipd,    WRDATA2,        tipd_WRDATA2);
        VitalWireDelay (WRDATA3_ipd,    WRDATA3,        tipd_WRDATA3);
        VitalWireDelay (RAD0_ipd,              RAD0,          tipd_RAD0);
        VitalWireDelay (RAD1_ipd,              RAD1,          tipd_RAD1);
        VitalWireDelay (RAD2_ipd,              RAD2,          tipd_RAD2);
        VitalWireDelay (RAD3_ipd,              RAD3,          tipd_RAD3);
        VitalWireDelay (RAD4_ipd,              RAD4,          tipd_RAD4);
        VitalWireDelay (WRAD0_ipd,              WRAD0,          tipd_WRAD0);
        VitalWireDelay (WRAD1_ipd,              WRAD1,          tipd_WRAD1);
        VitalWireDelay (WRAD2_ipd,              WRAD2,          tipd_WRAD2);
        VitalWireDelay (WRAD3_ipd,              WRAD3,          tipd_WRAD3);
        VitalWireDelay (WRAD4_ipd,              WRAD4,          tipd_WRAD4);
  END BLOCK;

  ---------------------------------------------------------------------
  -- Behavior Section
  ---------------------------------------------------------------------

  ---------------------------------------------------------------------
  -- Wrapper Section
  ---------------------------------------------------------------------

   wrapper_read_add : process(REN_ipd, RAD4_ipd, RAD3_ipd, RAD2_ipd, RAD1_ipd, RAD0_ipd, WEN_ipd)

   begin
    if (REN_ipd = '1') then
        RD_ADD(4) <= RAD4_ipd;
        RD_ADD(3) <= RAD3_ipd;
        RD_ADD(2) <= RAD2_ipd;
        RD_ADD(1) <= RAD1_ipd;
        RD_ADD(0) <= RAD0_ipd;
    else
	RD_ADD <= x_add;
    end if;

   end process;

   wrapper_read_add_w : process(REN_ipd, OE_ipd, WRAD4_ipd, WRAD3_ipd, WRAD2_ipd, WRAD1_ipd, WRAD0_ipd, WEN_ipd)

   begin
    if (REN_ipd = '1' and OE_ipd = '1' and WEN_ipd = '0') then
        RD_ADD_W(4) <= WRAD4_ipd;
        RD_ADD_W(3) <= WRAD3_ipd;
        RD_ADD_W(2) <= WRAD2_ipd;
        RD_ADD_W(1) <= WRAD1_ipd;
        RD_ADD_W(0) <= WRAD0_ipd;
    else
	RD_ADD_W <= x_add;
    end if;

   end process;

   wrapper_read_clk : process(REN_ipd, RCLK_ipd, WEN_ipd)

   begin
    if (REN_ipd = '1') then
	RD_CLK <= RCLK_ipd;
    else
	RD_CLK <= '0';
    end if;

   end process;

   wrapper_read_clk_w : process(REN_ipd, OE_ipd, WRCLK_ipd, WEN_ipd)

   begin
    if (REN_ipd = '1' and OE_ipd = '1' and WEN_ipd = '0') then
	RD_CLK_W <= WRCLK_ipd;
    else
	RD_CLK_W <= '0';
    end if;

   end process;

   wrapper_write_add : process(WEN_ipd, WRAD4_ipd, WRAD3_ipd, WRAD2_ipd, WRAD1_ipd, WRAD0_ipd)

   begin
    if (WEN_ipd = '1') then
        WR_ADD(4) <= WRAD4_ipd;
        WR_ADD(3) <= WRAD3_ipd;
        WR_ADD(2) <= WRAD2_ipd;
        WR_ADD(1) <= WRAD1_ipd;
        WR_ADD(0) <= WRAD0_ipd;
    else
	WR_ADD <= x_add;
    end if;

   end process;

   wrapper_write_clk : process(WEN_ipd, WRCLK_ipd)

   begin
    if (WEN_ipd = '1') then
	WR_CLK <= WRCLK_ipd;
    else
	WR_CLK <= '0';
    end if;

   end process;

   process(WR_CLK)

    begin
      if WR_CLK = '1' then
        write_add(4) <= WRAD4_ipd;
        write_add(3) <= WRAD3_ipd;
        write_add(2) <= WRAD2_ipd;
        write_add(1) <= WRAD1_ipd;
        write_add(0) <= WRAD0_ipd;
      end if;

   end process;

   wrapper_write_data : process(WEN_ipd, WRDATA3_ipd, WRDATA2_ipd, WRDATA1_ipd, WRDATA0_ipd)

   begin
    if (WEN_ipd = '1') then
        DIN(3) <= WRDATA3_ipd;
        DIN(2) <= WRDATA2_ipd;
        DIN(1) <= WRDATA1_ipd;
        DIN(0) <= WRDATA0_ipd;
    else
	DIN <= x_data;
    end if;

   end process;


  VITALBehavior : PROCESS ( WEN_ipd, REN_ipd, WR_CLK, RD_CLK_W, RD_CLK, DIN, RD_ADD, RD_ADD_W, WR_ADD )

   VARIABLE memory_array : memory_array_typ;
--   VARIABLE array_data_out : data_word_typ := x_data;
--   VARIABLE array_data_out_w : data_word_typ := z_data;

   -- Temporary variables
   VARIABLE tempaddr : integer := 0;
   VARIABLE rd_address : integer := 0;
   VARIABLE rd_address_w : integer := 0;

   -- Timing Check results
   VARIABLE Pviol_RCLK				: std_logic := '0';
   VARIABLE PeriodData_RCLK			: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_WRCLK				: std_logic := '0';
   VARIABLE PeriodData_WRCLK			: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_WR_ADD_stp_hld_0		: std_logic := '0';
   VARIABLE TimingData_WR_ADD_stp_hld_0		: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_WR_ADD_stp_hld_1		: std_logic := '0';
   VARIABLE TimingData_WR_ADD_stp_hld_1		: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_WR_ADD_stp_hld_2		: std_logic := '0';
   VARIABLE TimingData_WR_ADD_stp_hld_2		: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_WR_ADD_stp_hld_3		: std_logic := '0';
   VARIABLE TimingData_WR_ADD_stp_hld_3		: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_WR_ADD_stp_hld_4		: std_logic := '0';
   VARIABLE TimingData_WR_ADD_stp_hld_4		: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_WR_DATA_stp_0			: std_logic := '0';
   VARIABLE TimingData_WR_DATA_stp_0		: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_WR_DATA_stp_1			: std_logic := '0';
   VARIABLE TimingData_WR_DATA_stp_1		: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_WR_DATA_stp_2			: std_logic := '0';
   VARIABLE TimingData_WR_DATA_stp_2		: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_WR_DATA_stp_3			: std_logic := '0';
   VARIABLE TimingData_WR_DATA_stp_3		: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_WR_DATA_hld_0			: std_logic := '0';
   VARIABLE TimingData_WR_DATA_hld_0		: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_WR_DATA_hld_1			: std_logic := '0';
   VARIABLE TimingData_WR_DATA_hld_1		: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_WR_DATA_hld_2			: std_logic := '0';
   VARIABLE TimingData_WR_DATA_hld_2		: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_WR_DATA_hld_3			: std_logic := '0';
   VARIABLE TimingData_WR_DATA_hld_3		: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_RD_ADD_stp_hld_0		: std_logic := '0';
   VARIABLE TimingData_RD_ADD_stp_hld_0		: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_RD_ADD_stp_hld_1		: std_logic := '0';
   VARIABLE TimingData_RD_ADD_stp_hld_1		: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_RD_ADD_stp_hld_2		: std_logic := '0';
   VARIABLE TimingData_RD_ADD_stp_hld_2		: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_RD_ADD_stp_hld_3		: std_logic := '0';
   VARIABLE TimingData_RD_ADD_stp_hld_3		: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_RD_ADD_stp_hld_4		: std_logic := '0';
   VARIABLE TimingData_RD_ADD_stp_hld_4		: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_WEN_hld			: std_logic := '0';
   VARIABLE TimingData_WEN_hld			: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_REN_hld			: std_logic := '0';
   VARIABLE TimingData_REN_hld			: VitalTimingDataType := VitalTimingDataInit;



 BEGIN

    -- Timing Check Section
    -------------------------------------------------------------------
    IF (TimingChecksOn) THEN

        VitalSetupHoldCheck    (Tviol_WR_ADD_stp_hld_0,
                                TimingData_WR_ADD_stp_hld_0,
                                WR_ADD(0), "WRAD0",
                                0.0 ns,
                                WR_CLK, "WRCLK",
                                0.0 ns,
                                tsetup_WRAD0_WRCLK_noedge_posedge, tsetup_WRAD0_WRCLK_noedge_posedge,
                                thold_WRAD0_WRCLK_noedge_posedge, thold_WRAD0_WRCLK_noedge_posedge,
                                WEN_ipd = '1',
                                '/',
                                InstancePath & "/RB_DS",
                                TRUE,
                                TRUE,
                                WARNING );

        VitalSetupHoldCheck    (Tviol_WR_ADD_stp_hld_1,
                                TimingData_WR_ADD_stp_hld_1,
                                WR_ADD(1), "WRAD1",
                                0.0 ns,
                                WR_CLK, "WRCLK",
                                0.0 ns,
                                tsetup_WRAD1_WRCLK_noedge_posedge, tsetup_WRAD1_WRCLK_noedge_posedge,
                                thold_WRAD1_WRCLK_noedge_posedge, thold_WRAD1_WRCLK_noedge_posedge,
                                WEN_ipd = '1',
                                '/',
                                InstancePath & "/RB_DS",
                                TRUE,
                                TRUE,
                                WARNING );

        VitalSetupHoldCheck    (Tviol_WR_ADD_stp_hld_2,
                                TimingData_WR_ADD_stp_hld_2,
                                WR_ADD(2), "WRAD2",
                                0.0 ns,
                                WR_CLK, "WRCLK",
                                0.0 ns,
                                tsetup_WRAD2_WRCLK_noedge_posedge, tsetup_WRAD2_WRCLK_noedge_posedge,
                                thold_WRAD2_WRCLK_noedge_posedge, thold_WRAD2_WRCLK_noedge_posedge,
                                WEN_ipd = '1',
                                '/',
                                InstancePath & "/RB_DS",
                                TRUE,
                                TRUE,
                                WARNING );
       VitalSetupHoldCheck    (Tviol_WR_ADD_stp_hld_3,
                                TimingData_WR_ADD_stp_hld_3,
                                WR_ADD(3), "WRAD3",
                                0.0 ns,
                                WR_CLK, "WRCLK",
                                0.0 ns,
                                tsetup_WRAD3_WRCLK_noedge_posedge, tsetup_WRAD3_WRCLK_noedge_posedge,
                                thold_WRAD3_WRCLK_noedge_posedge, thold_WRAD3_WRCLK_noedge_posedge,
                                WEN_ipd = '1',
                                '/',
                                InstancePath & "/RB_DS",
                                TRUE,
                                TRUE,
                                WARNING );
        VitalSetupHoldCheck    (Tviol_WR_ADD_stp_hld_4,
                                TimingData_WR_ADD_stp_hld_4,
                                WR_ADD(4), "WRAD4",
                                0.0 ns,
                                WR_CLK, "WRCLK",
                                0.0 ns,
                                tsetup_WRAD4_WRCLK_noedge_posedge, tsetup_WRAD4_WRCLK_noedge_posedge,
                                thold_WRAD4_WRCLK_noedge_posedge, thold_WRAD4_WRCLK_noedge_posedge,
                                WEN_ipd = '1',
                                '/',
                                InstancePath & "/RB_DS",
                                TRUE,
                                TRUE,
                                WARNING );

        VitalSetupHoldCheck    (Tviol_WR_DATA_stp_0,
                                TimingData_WR_DATA_stp_0,
                                DIN(0), "WRDATA0",
                                0.0 ns,
                                WR_CLK, "WRCLK",
                                0.0 ns,
                                tsetup_WRDATA0_WRCLK_noedge_posedge, tsetup_WRDATA0_WRCLK_noedge_posedge,
                                0.0 ns, 0.0 ns,
                                WEN_ipd = '1',
                                '/',
                                InstancePath & "/RB_DS",
                                TRUE,
                                TRUE,
                                WARNING );

        VitalSetupHoldCheck    (Tviol_WR_DATA_stp_1,
                                TimingData_WR_DATA_stp_1,
                                DIN(1), "WRDATA1",
                                0.0 ns,
                                WR_CLK, "WRCLK",
                                0.0 ns,
                                tsetup_WRDATA1_WRCLK_noedge_posedge, tsetup_WRDATA1_WRCLK_noedge_posedge,
                                0.0 ns, 0.0 ns,
                                WEN_ipd = '1',
                                '/',
                                InstancePath & "/RB_DS",
                                TRUE,
                                TRUE,
                                WARNING );

        VitalSetupHoldCheck    (Tviol_WR_DATA_stp_2,
                                TimingData_WR_DATA_stp_2,
                                DIN(2), "WRDATA2",
                                0.0 ns,
                                WR_CLK, "WRCLK",
                                0.0 ns,
                                tsetup_WRDATA2_WRCLK_noedge_posedge, tsetup_WRDATA2_WRCLK_noedge_posedge,
                                0.0 ns, 0.0 ns,
                                WEN_ipd = '1',
                                '/',
                                InstancePath & "/RB_DS",
                                TRUE,
                                TRUE,
                                WARNING );
       VitalSetupHoldCheck    (Tviol_WR_DATA_stp_3,
                                TimingData_WR_DATA_stp_3,
                                DIN(3), "WRDATA3",
                                0.0 ns,
                                WR_CLK, "WRCLK",
                                0.0 ns,
                                tsetup_WRDATA3_WRCLK_noedge_posedge, tsetup_WRDATA3_WRCLK_noedge_posedge,
                                0.0 ns, 0.0 ns,
                                WEN_ipd = '1',
                                '/',
                                InstancePath & "/RB_DS",
                                TRUE,
                                TRUE,
                                WARNING );

        VitalSetupHoldCheck    (Tviol_WR_DATA_hld_0,
                                TimingData_WR_DATA_hld_0,
                                DIN(0), "WRDATA0",
                                0.0 ns,
                                WR_CLK, "WRCLK",
                                0.0 ns,
                                0.0 ns, 0.0 ns,
                                thold_WRDATA0_WRCLK_noedge_posedge, thold_WRDATA0_WRCLK_noedge_posedge,
                                WEN_ipd = '1',
                                '/',
                                InstancePath & "/RB_DS",
                                TRUE,
                                TRUE,
                                WARNING );

        VitalSetupHoldCheck    (Tviol_WR_DATA_hld_1,
                                TimingData_WR_DATA_hld_1,
                                DIN(1), "WRDATA1",
                                0.0 ns,
                                WR_CLK, "WRCLK",
                                0.0 ns,
                                0.0 ns, 0.0 ns,
                                thold_WRDATA1_WRCLK_noedge_posedge, thold_WRDATA1_WRCLK_noedge_posedge,
                                WEN_ipd = '1',
                                '/',
                                InstancePath & "/RB_DS",
                                TRUE,
                                TRUE,
                                WARNING );

        VitalSetupHoldCheck    (Tviol_WR_DATA_hld_2,
                                TimingData_WR_DATA_hld_2,
                                DIN(2), "WRDATA2",
                                0.0 ns,
                                WR_CLK, "WRCLK",
                                0.0 ns,
                                0.0 ns, 0.0 ns,
                                thold_WRDATA2_WRCLK_noedge_posedge, thold_WRDATA2_WRCLK_noedge_posedge,
                                WEN_ipd = '1',
                                '/',
                                InstancePath & "/RB_DS",
                                TRUE,
                                TRUE,
                                WARNING );
        VitalSetupHoldCheck    (Tviol_WR_DATA_hld_3,
                                TimingData_WR_DATA_hld_3,
                                DIN(3), "WRDATA3",
                                0.0 ns,
                                WR_CLK, "WRCLK",
                                0.0 ns,
                                0.0 ns, 0.0 ns,
                                thold_WRDATA3_WRCLK_noedge_posedge, thold_WRDATA3_WRCLK_noedge_posedge,
                                WEN_ipd = '1',
                                '/',
                                InstancePath & "/RB_DS",
                                TRUE,
                                TRUE,
                                WARNING );


        VitalSetupHoldCheck    (Tviol_WEN_hld,
                                TimingData_WEN_hld,
                                WEN_ipd, "WEN",
                                0.0 ns,
                                WR_CLK, "WRCLK",
                                0.0 ns,
                                tsetup_WEN_WRCLK_noedge_posedge, tsetup_WEN_WRCLK_noedge_posedge,
                                thold_WEN_WRCLK_noedge_posedge, thold_WEN_WRCLK_noedge_posedge,
                                True,
                                '/',
                                InstancePath & "/RB_DS",
                                TRUE,
                                TRUE,
                                WARNING );

	VitalPeriodPulseCheck  (Pviol_RCLK,
				PeriodData_RCLK,
				RCLK_ipd, "RCLK",
				0.0 ns,
				0.0 ns,
				tpw_RCLK_posedge,
				0.0 ns,
				TRUE,
				InstancePath & "/RB_DS",
				TRUE,
				TRUE,
				WARNING );

	VitalPeriodPulseCheck  (Pviol_WRCLK,
				PeriodData_WRCLK,
				WRCLK_ipd, "WRCLK",
				0.0 ns,
				0.0 ns,
				tpw_WRCLK_posedge,
				0.0 ns,
				TRUE,
				InstancePath & "/RB_DS",
				TRUE,
				TRUE,
				WARNING );


        VitalSetupHoldCheck    (Tviol_RD_ADD_stp_hld_0,
                                TimingData_RD_ADD_stp_hld_0,
                                RD_ADD(0), "RAD0",
                                0.0 ns,
                                RD_CLK, "RCLK",
                                0.0 ns,
                                tsetup_RAD0_RCLK_noedge_posedge, tsetup_RAD0_RCLK_noedge_posedge,
                                thold_RAD0_RCLK_noedge_posedge, thold_RAD0_RCLK_noedge_posedge,
                                REN_ipd = '1' ,
                                '/',
                                InstancePath & "/RB_DS",
                                TRUE,
                                TRUE,
                                WARNING );

        VitalSetupHoldCheck    (Tviol_RD_ADD_stp_hld_1,
                                TimingData_RD_ADD_stp_hld_1,
                                RD_ADD(1), "RAD1",
                                0.0 ns,
                                RD_CLK, "RCLK",
                                0.0 ns,
                                tsetup_RAD1_RCLK_noedge_posedge, tsetup_RAD1_RCLK_noedge_posedge,
                                thold_RAD1_RCLK_noedge_posedge, thold_RAD1_RCLK_noedge_posedge,
                                REN_ipd = '1' ,
                                '/',
                                InstancePath & "/RB_DS",
                                TRUE,
                                TRUE,
                                WARNING );

        VitalSetupHoldCheck    (Tviol_RD_ADD_stp_hld_2,
                                TimingData_RD_ADD_stp_hld_2,
                                RD_ADD(2), "RAD2",
                                0.0 ns,
                                RD_CLK, "RCLK",
                                0.0 ns,
                                tsetup_RAD2_RCLK_noedge_posedge, tsetup_RAD2_RCLK_noedge_posedge,
                                thold_RAD2_RCLK_noedge_posedge, thold_RAD2_RCLK_noedge_posedge,
                                REN_ipd = '1' ,
                                '/',
                                InstancePath & "/RB_DS",
                                TRUE,
                                TRUE,
                                WARNING );

        VitalSetupHoldCheck    (Tviol_RD_ADD_stp_hld_3,
                                TimingData_RD_ADD_stp_hld_3,
                                RD_ADD(3), "RAD3",
                                0.0 ns,
                                RD_CLK, "RCLK",
                                0.0 ns,
                                tsetup_RAD3_RCLK_noedge_posedge, tsetup_RAD3_RCLK_noedge_posedge,
                                thold_RAD3_RCLK_noedge_posedge, thold_RAD3_RCLK_noedge_posedge,
                                REN_ipd = '1' ,
                                '/',
                                InstancePath & "/RB_DS",
                                TRUE,
                                TRUE,
                                WARNING );
        VitalSetupHoldCheck    (Tviol_RD_ADD_stp_hld_4,
                                TimingData_RD_ADD_stp_hld_4,
                                RD_ADD(4), "RAD4",
                                0.0 ns,
                                RD_CLK, "RCLK",
                                0.0 ns,
                                tsetup_RAD4_RCLK_noedge_posedge, tsetup_RAD4_RCLK_noedge_posedge,
                                thold_RAD4_RCLK_noedge_posedge, thold_RAD4_RCLK_noedge_posedge,
                                REN_ipd = '1' ,
                                '/',
                                InstancePath & "/RB_DS",
                                TRUE,
                                TRUE,
                                WARNING );

        VitalSetupHoldCheck    (Tviol_REN_hld,
                                TimingData_REN_hld,
                                REN_ipd, "REN",
                                0.0 ns,
                                RD_CLK, "RCLK",
                                0.0 ns,
                                tsetup_REN_RCLK_noedge_posedge, tsetup_REN_RCLK_noedge_posedge,
                                thold_REN_RCLK_noedge_posedge, thold_REN_RCLK_noedge_posedge,
                                True,
                                '/',
                                InstancePath & "/RB_DS",
                                TRUE,
                                TRUE,
                                WARNING );


    END IF; -- Timing Check Section

    -------------------------------------------------------------------
    -- Functionality Section
    -------------------------------------------------------------------

-- WRITE ADDRESS GOES XX

    if ( WR_CLK'EVENT and WR_CLK = '1' and vecX(WR_ADD)) then

        assert false
        report "Illegal Address Input: Undefined  Address at the Read_Write Port."
        severity note ;
        memory_array := (others => x_data);

    end if;

-- ADDRESS HOLD AND SETUP VIOLATION EFFECT

    if( Tviol_WR_ADD_stp_hld_0 = 'X' or Tviol_WR_ADD_stp_hld_1 = 'X' or Tviol_WR_ADD_stp_hld_2 = 'X' or Tviol_WR_ADD_stp_hld_3 = 'X' or Tviol_WR_ADD_stp_hld_4 = 'X' ) then
	memory_array := (others => x_data);
    else
 
-- DATA SETUP AND HOLD VIOLATION EFFECT

    if( Pviol_WRCLK = 'X' or Tviol_WR_DATA_hld_0 = 'X' or Tviol_WR_DATA_hld_1 = 'X' or Tviol_WR_DATA_hld_2 = 'X' or Tviol_WR_DATA_hld_3 = 'X' or Tviol_WEN_hld = 'X') then
	tempaddr := vec2int(write_add);
	memory_array(tempaddr) := x_data;
    end if;

    if( Tviol_WR_DATA_stp_0 = 'X' or Tviol_WR_DATA_stp_1 = 'X' or Tviol_WR_DATA_stp_2 = 'X' or Tviol_WR_DATA_stp_3 = 'X') then
	tempaddr := vec2int(WR_ADD);
	memory_array(tempaddr) := x_data;
    end if;

    end if;

-- VALID MEMORY WRITE

    if ( WR_CLK'EVENT and WR_CLK = '1' and not vecX(WR_ADD) and not( Tviol_WR_ADD_stp_hld_0 = 'X' or Tviol_WR_ADD_stp_hld_1 = 'X' or Tviol_WR_ADD_stp_hld_2 = 'X' or Tviol_WR_ADD_stp_hld_3 = 'X' or Tviol_WR_ADD_stp_hld_4 = 'X' ) and not ( Pviol_WRCLK = 'X' or Tviol_WR_DATA_hld_0 = 'X' or Tviol_WR_DATA_hld_1 = 'X' or Tviol_WR_DATA_hld_2 = 'X' or Tviol_WR_DATA_hld_3 = 'X' or Tviol_WEN_hld = 'X') and not( Tviol_WR_DATA_stp_0 = 'X' or Tviol_WR_DATA_stp_1 = 'X' or Tviol_WR_DATA_stp_2 = 'X' or Tviol_WR_DATA_stp_3 = 'X') ) then
	tempaddr := vec2int(WR_ADD);
	memory_array(tempaddr) := DIN;
    end if;

    if WR_CLK'EVENT and WR_CLK /= WRCLK_ipd and WR_CLK'LAST_VALUE = '1' then
	memory_array(tempaddr) := x_data;
    end if;


-- READ ADDRESS CYCLE VIOLATION EFFECT

    if( Tviol_RD_ADD_stp_hld_0 = 'X' or Tviol_RD_ADD_stp_hld_1 = 'X' or Tviol_RD_ADD_stp_hld_2 = 'X' or Tviol_RD_ADD_stp_hld_3 = 'X' or Tviol_RD_ADD_stp_hld_4 = 'X' or Pviol_RCLK = 'X' or Tviol_REN_hld = 'X' or (RD_CLK'EVENT and RD_CLK = '1' and vecX(RD_ADD))) then
	data_out <= x_data;
    elsif


-- VALID MEMORY READ

    (RD_CLK'EVENT and RD_CLK = '1' and not( Tviol_RD_ADD_stp_hld_0 = 'X' or Tviol_RD_ADD_stp_hld_1 = 'X' or Tviol_RD_ADD_stp_hld_2 = 'X' or Tviol_RD_ADD_stp_hld_3 = 'X' or Tviol_RD_ADD_stp_hld_4 = 'X' or Pviol_RCLK = 'X' or Tviol_REN_hld = 'X' or vecX(RD_ADD) )) then
	rd_address := vec2int(RD_ADD);
	data_out <= memory_array(rd_address);
    end if;

    if RD_CLK'EVENT and RD_CLK /= RCLK_ipd and RD_CLK'LAST_VALUE = '1' then
	data_out <= x_data;
    end if;


-- READ ADDRESS CYCLE VIOLATION EFFECT

    if( Tviol_WR_ADD_stp_hld_0 = 'X' or Tviol_WR_ADD_stp_hld_1 = 'X' or Tviol_WR_ADD_stp_hld_2 = 'X' or Tviol_WR_ADD_stp_hld_3 = 'X' or Tviol_WR_ADD_stp_hld_4 = 'X' or Pviol_WRCLK = 'X' or Tviol_REN_hld  = 'X' or (RD_CLK_W'EVENT and RD_CLK_W = '1' and vecX(RD_ADD_W)) ) then
	data_out_w <= x_data;
    elsif

-- VALID MEMORY READ

    (RD_CLK_W'EVENT and RD_CLK_W = '1' and not( Tviol_WR_ADD_stp_hld_0 = 'X' or Tviol_WR_ADD_stp_hld_1 = 'X' or Tviol_WR_ADD_stp_hld_2 = 'X' or Tviol_WR_ADD_stp_hld_3 = 'X' or Tviol_WR_ADD_stp_hld_4 = 'X' or Pviol_WRCLK = 'X' or Tviol_REN_hld = 'X' or vecX(RD_ADD_W) ))then
	rd_address_w := vec2int(RD_ADD_W);
	data_out_w <= memory_array(rd_address_w);
    end if;

    if RD_CLK_W'EVENT and RD_CLK_W /= WRCLK_ipd and RD_CLK_W'LAST_VALUE = '1' then
	data_out_w <= x_data;
    end if;

--data_out <= array_data_out;

--data_out_w <= array_data_out_w;


  END PROCESS;

    -------------------------------------------------------------------------------
    -- Temporary output signal should get assigned to the output signal.
    -------------------------------------------------------------------------------

PROCESS(data_out_w, WRCLK_ipd, OE_ipd)

   VARIABLE GLITCH_DATA : VitalGlitchDataType;
   VARIABLE con : std_logic ;--:= '0';
    VARIABLE WEN_inv : std_logic ;--:= '0';
    VARIABLE WRDATA3_1 : std_logic := 'Z';
    VARIABLE WRDATA2_1 : std_logic := 'Z';
    VARIABLE WRDATA1_1 : std_logic := 'Z';
    VARIABLE WRDATA0_1 : std_logic := 'Z';

   BEGIN
       WEN_inv := VitalINV(WEN_ipd);
       con := VitalAND3(OE_ipd,REN_ipd, WEN_inv);


      WRDATA3_1 := VITALBUFIF1(data_out_w(3),con);
      WRDATA2_1 := VITALBUFIF1(data_out_w(2),con);
      WRDATA1_1 := VITALBUFIF1(data_out_w(1),con);
      WRDATA0_1 := VITALBUFIF1(data_out_w(0),con);


      VitalPathDelay01Z ( WRDATA0, GLITCH_DATA, "WRDATA0", WRDATA0_1,
        Paths => (
        0 => ( WRCLK_ipd'LAST_EVENT, tpd_WRCLK_WRDATA0, TRUE),
        1 => ( OE_ipd'LAST_EVENT, tpd_OE_WRDATA0, TRUE )),
        DefaultDelay=>VitalZeroDelay01Z,
        Mode=>VitalInertial,
        XON=>TRUE,
        MsgOn=>TRUE,
        MsgSeverity=>WARNING );

      VitalPathDelay01Z ( WRDATA1, GLITCH_DATA, "WRDATA1", WRDATA1_1,
        Paths => (
        0 => ( WRCLK_ipd'LAST_EVENT, tpd_WRCLK_WRDATA1, TRUE),
        1 => ( OE_ipd'LAST_EVENT, tpd_OE_WRDATA1, TRUE )),
        DefaultDelay=>VitalZeroDelay01Z,
        Mode=>VitalInertial,
        XON=>TRUE,
        MsgOn=>TRUE,
        MsgSeverity=>WARNING );

      VitalPathDelay01Z ( WRDATA2, GLITCH_DATA, "WRDATA2", WRDATA2_1,
        Paths => (
        0 => ( WRCLK_ipd'LAST_EVENT, tpd_WRCLK_WRDATA2, TRUE),
        1 => ( OE_ipd'LAST_EVENT, tpd_OE_WRDATA2, TRUE )),
        DefaultDelay=>VitalZeroDelay01Z,
        Mode=>VitalInertial,
        XON=>TRUE,
        MsgOn=>TRUE,
        MsgSeverity=>WARNING );

      VitalPathDelay01Z ( WRDATA3, GLITCH_DATA, "WRDATA3", WRDATA3_1,
        Paths => (
        0 => ( WRCLK_ipd'LAST_EVENT, tpd_WRCLK_WRDATA3, TRUE),
        1 => ( OE_ipd'LAST_EVENT, tpd_OE_WRDATA3, TRUE )),
        DefaultDelay=>VitalZeroDelay01Z,
        Mode=>VitalInertial,
        XON=>TRUE,
        MsgOn=>TRUE,
        MsgSeverity=>WARNING );

END PROCESS;

PROCESS(data_out, RCLK_ipd)

    VARIABLE RDATA3_1 : std_logic := 'X';--:= 'X';
    VARIABLE RDATA2_1 : std_logic := 'X';--:= 'X';
    VARIABLE RDATA1_1 : std_logic := 'X';--:= 'X';
    VARIABLE RDATA0_1 : std_logic := 'X';--:= 'X';
    VARIABLE GLITCH : VitalGlitchDataType;
    BEGIN

      RDATA3_1 := VITALBUF(data_out(3));
      RDATA2_1 := VITALBUF(data_out(2));
      RDATA1_1 := VITALBUF(data_out(1));
      RDATA0_1 := VITALBUF(data_out(0));

      VitalPathDelay01 ( RDATA3, GLITCH, "RDATA3", RDATA3_1,
        Paths => (
        0 => ( RCLK_ipd'LAST_EVENT, tpd_RCLK_RDATA3, TRUE )),
        DefaultDelay=>VitalZeroDelay01,
        Mode=>VitalInertial,
        XON=>TRUE,
        MsgOn=>TRUE,
        MsgSeverity=>WARNING );

      VitalPathDelay01 ( RDATA2, GLITCH, "RDATA2", RDATA2_1,
        Paths => (
        0 => ( RCLK_ipd'LAST_EVENT, tpd_RCLK_RDATA2, TRUE )),
        DefaultDelay=>VitalZeroDelay01,
        Mode=>VitalInertial,
        XON=>TRUE,
        MsgOn=>TRUE,
        MsgSeverity=>WARNING );

      VitalPathDelay01 ( RDATA1, GLITCH, "RDATA1", RDATA1_1,
        Paths => (
        0 => ( RCLK_ipd'LAST_EVENT, tpd_RCLK_RDATA1, TRUE )),
        DefaultDelay=>VitalZeroDelay01,
        Mode=>VitalInertial,
        XON=>TRUE,
        MsgOn=>TRUE,
        MsgSeverity=>WARNING );

      VitalPathDelay01 ( RDATA0, GLITCH, "RDATA0", RDATA0_1,
        Paths => (
        0 => ( RCLK_ipd'LAST_EVENT, tpd_RCLK_RDATA0, TRUE )),
        DefaultDelay=>VitalZeroDelay01,
        Mode=>VitalInertial,
        XON=>TRUE,
        MsgOn=>TRUE,
        MsgSeverity=>WARNING );

END PROCESS;

END VITAL_VF;
configuration CFG_RB_DS_VITAL of RB_DS is
        for VITAL_VF
        end for;
end CFG_RB_DS_VITAL;
-----------------------------------------------------------------------

-- VITAL model for RB_MA 30.10 technology
-----------------------------------------------------------------------

LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.VITAL_timing.all;
USE IEEE.VITAL_primitives.all;
LIBRARY VF1;
USE VF1.ALL;
USE VF1.RAMPACK.ALL;

-----------------------------------------------------------------------
-- ENTITY declaration
-----------------------------------------------------------------------

ENTITY RB_MA IS
  GENERIC (
	tipd_WEN		: VitalDelayType01			:= (0.0 ns, 0.0 ns);
	tipd_WRCLK		: VitalDelayType01			:= (0.0 ns, 0.0 ns);
	tipd_OE		: VitalDelayType01			:= (0.0 ns, 0.0 ns);
        tipd_WRDATA3            : VitalDelayType01      := (0.0 ns, 0.0 ns);
        tipd_WRDATA2            : VitalDelayType01      := (0.0 ns, 0.0 ns);
        tipd_WRDATA1            : VitalDelayType01      := (0.0 ns, 0.0 ns);
        tipd_WRDATA0            : VitalDelayType01      := (0.0 ns, 0.0 ns);
        tipd_WRAD4              : VitalDelayType01      := (0.0 ns, 0.0 ns);
        tipd_WRAD3              : VitalDelayType01      := (0.0 ns, 0.0 ns);
        tipd_WRAD2              : VitalDelayType01      := (0.0 ns, 0.0 ns);
        tipd_WRAD1              : VitalDelayType01      := (0.0 ns, 0.0 ns);
        tipd_WRAD0              : VitalDelayType01      := (0.0 ns, 0.0 ns);

tpw_WRCLK_posedge        :VitalDelayType := 1.0 ns;
tsetup_WRDATA3_WRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
thold_WRDATA3_WRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
tsetup_WRDATA2_WRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
thold_WRDATA2_WRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
tsetup_WRDATA1_WRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
thold_WRDATA1_WRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
tsetup_WRDATA0_WRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
thold_WRDATA0_WRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
tsetup_WRAD4_WRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
thold_WRAD4_WRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
tsetup_WRAD3_WRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
thold_WRAD3_WRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
tsetup_WRAD2_WRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
thold_WRAD2_WRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
tsetup_WRAD1_WRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
thold_WRAD1_WRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
tsetup_WRAD0_WRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
thold_WRAD0_WRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
tsetup_WEN_WRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
thold_WEN_WRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;

tpd_WRAD4_WRDATA0         :VitalDelayType01Z := (2 ns,2 ns,2 ns,2 ns,2 ns,2 ns);
tpd_WRAD3_WRDATA0         :VitalDelayType01Z := (2 ns,2 ns,2 ns,2 ns,2 ns,2 ns);
tpd_WRAD2_WRDATA0         :VitalDelayType01Z := (2 ns,2 ns,2 ns,2 ns,2 ns,2 ns);
tpd_WRAD1_WRDATA0         :VitalDelayType01Z := (2 ns,2 ns,2 ns,2 ns,2 ns,2 ns);
tpd_WRAD0_WRDATA0         :VitalDelayType01Z := (2 ns,2 ns,2 ns,2 ns,2 ns,2 ns);
tpd_WRAD4_WRDATA1         :VitalDelayType01Z := (2 ns,2 ns,2 ns,2 ns,2 ns,2 ns);
tpd_WRAD3_WRDATA1         :VitalDelayType01Z := (2 ns,2 ns,2 ns,2 ns,2 ns,2 ns);
tpd_WRAD2_WRDATA1         :VitalDelayType01Z := (2 ns,2 ns,2 ns,2 ns,2 ns,2 ns);
tpd_WRAD1_WRDATA1         :VitalDelayType01Z := (2 ns,2 ns,2 ns,2 ns,2 ns,2 ns);
tpd_WRAD0_WRDATA1         :VitalDelayType01Z := (2 ns,2 ns,2 ns,2 ns,2 ns,2 ns);
tpd_WRAD4_WRDATA2         :VitalDelayType01Z := (2 ns,2 ns,2 ns,2 ns,2 ns,2 ns);
tpd_WRAD3_WRDATA2         :VitalDelayType01Z := (2 ns,2 ns,2 ns,2 ns,2 ns,2 ns);
tpd_WRAD2_WRDATA2         :VitalDelayType01Z := (2 ns,2 ns,2 ns,2 ns,2 ns,2 ns);
tpd_WRAD1_WRDATA2         :VitalDelayType01Z := (2 ns,2 ns,2 ns,2 ns,2 ns,2 ns);
tpd_WRAD0_WRDATA2         :VitalDelayType01Z := (2 ns,2 ns,2 ns,2 ns,2 ns,2 ns);
tpd_WRAD4_WRDATA3         :VitalDelayType01Z := (2 ns,2 ns,2 ns,2 ns,2 ns,2 ns);
tpd_WRAD3_WRDATA3         :VitalDelayType01Z := (2 ns,2 ns,2 ns,2 ns,2 ns,2 ns);
tpd_WRAD2_WRDATA3         :VitalDelayType01Z := (2 ns,2 ns,2 ns,2 ns,2 ns,2 ns);
tpd_WRAD1_WRDATA3         :VitalDelayType01Z := (2 ns,2 ns,2 ns,2 ns,2 ns,2 ns);
tpd_WRAD0_WRDATA3         :VitalDelayType01Z := (2 ns,2 ns,2 ns,2 ns,2 ns,2 ns);
tpd_OE_WRDATA0         :VitalDelayType01Z := (2 ns,2 ns,2 ns,2 ns,2 ns,2 ns);
tpd_OE_WRDATA1         :VitalDelayType01Z := (2 ns,2 ns,2 ns,2 ns,2 ns,2 ns);
tpd_OE_WRDATA2         :VitalDelayType01Z := (2 ns,2 ns,2 ns,2 ns,2 ns,2 ns);
tpd_OE_WRDATA3         :VitalDelayType01Z := (2 ns,2 ns,2 ns,2 ns,2 ns,2 ns);

	TimingChecksOn : BOOLEAN := TRUE;
	InstancePath : STRING := "*"
            );
  PORT	(
	WEN		: IN	std_logic ;
	WRCLK		: IN	std_logic ;
	OE		: IN	std_logic ;
        WRDATA3 : INOUT std_logic := 'Z';
        WRDATA2 : INOUT std_logic := 'Z';
        WRDATA1 : INOUT std_logic := 'Z';
        WRDATA0 : INOUT std_logic := 'Z';
        WRAD4           : IN    std_logic;
        WRAD3           : IN    std_logic;
        WRAD2           : IN    std_logic;
        WRAD1           : IN    std_logic;
        WRAD0           : IN    std_logic
	);


   ATTRIBUTE VITAL_LEVEL0 OF RB_MA : ENTITY IS TRUE;

END RB_MA;

-----------------------------------------------------------------------
-- ARCHITECTURE declaration
-----------------------------------------------------------------------
ARCHITECTURE VITAL_VF OF RB_MA IS

    ATTRIBUTE VITAL_LEVEL1 OF VITAL_VF : ARCHITECTURE IS FALSE;

	SIGNAL WEN_ipd		: std_logic := 'X';
	SIGNAL WRCLK_ipd		: std_logic := '0';
	SIGNAL WR_CLK		: std_logic := '0';
	SIGNAL OE_ipd	: std_logic := 'X';
	SIGNAL WR_ADD		: std_logic_vector(4 DOWNTO 0);
	SIGNAL write_add	: std_logic_vector(4 DOWNTO 0);
	SIGNAL data_out		: std_logic_vector(3 DOWNTO 0) := z_data;
	SIGNAL output_delay	: time		:= 0 ns;
        SIGNAL WRDATA3_ipd      : std_logic := 'Z';
        SIGNAL WRDATA2_ipd      : std_logic := 'Z';
        SIGNAL WRDATA1_ipd      : std_logic := 'Z';
        SIGNAL WRDATA0_ipd      : std_logic := 'Z';
        SIGNAL DIN              : std_logic_vector(3 DOWNTO 0);
        SIGNAL RD_ADD           : std_logic_vector(4 DOWNTO 0);
        SIGNAL WRAD4_ipd                : std_logic := '0';
        SIGNAL WRAD3_ipd                : std_logic := '0';
        SIGNAL WRAD2_ipd                : std_logic := '0';
        SIGNAL WRAD1_ipd                : std_logic := '0';
        SIGNAL WRAD0_ipd                : std_logic := '0';
	SIGNAL memory_array	: memory_array_typ;

BEGIN
   
  ---------------------------------------------------------------------
  -- INPUT PATH DELAYs
  ---------------------------------------------------------------------
  WIREDELAY : BLOCK
  BEGIN
	VitalWireDelay (WEN_ipd,		WEN,		tipd_WEN);
	VitalWireDelay (WRCLK_ipd,		WRCLK,		tipd_WRCLK);
	VitalWireDelay (OE_ipd,		OE,		tipd_OE);
        VitalWireDelay (WRDATA0_ipd,    WRDATA0,        tipd_WRDATA0);
        VitalWireDelay (WRDATA1_ipd,    WRDATA1,        tipd_WRDATA1);
        VitalWireDelay (WRDATA2_ipd,    WRDATA2,        tipd_WRDATA2);
        VitalWireDelay (WRDATA3_ipd,    WRDATA3,        tipd_WRDATA3);
        VitalWireDelay (WRAD0_ipd,              WRAD0,          tipd_WRAD0);
        VitalWireDelay (WRAD1_ipd,              WRAD1,          tipd_WRAD1);
        VitalWireDelay (WRAD2_ipd,              WRAD2,          tipd_WRAD2);
        VitalWireDelay (WRAD3_ipd,              WRAD3,          tipd_WRAD3);
        VitalWireDelay (WRAD4_ipd,              WRAD4,          tipd_WRAD4);

  END BLOCK;

  ---------------------------------------------------------------------
  -- Behavior Section
  ---------------------------------------------------------------------

  ---------------------------------------------------------------------
  -- Wrapper Section
  ---------------------------------------------------------------------

   wrapper_read_add : process(WEN_ipd, WRAD4_ipd, WRAD3_ipd, WRAD2_ipd, WRAD1_ipd, WRAD0_ipd)

   begin
    if (WEN_ipd = '0') then
        RD_ADD(4) <= WRAD4_ipd;
        RD_ADD(3) <= WRAD3_ipd;
        RD_ADD(2) <= WRAD2_ipd;
        RD_ADD(1) <= WRAD1_ipd;
        RD_ADD(0) <= WRAD0_ipd;
    else
	RD_ADD <= x_add;
    end if;

   end process;

   wrapper_write_add : process(WEN_ipd, WRAD4_ipd, WRAD3_ipd, WRAD2_ipd, WRAD1_ipd, WRAD0_ipd)

   begin
    if (WEN_ipd = '1') then
        WR_ADD(4) <= WRAD4_ipd;
        WR_ADD(3) <= WRAD3_ipd;
        WR_ADD(2) <= WRAD2_ipd;
        WR_ADD(1) <= WRAD1_ipd;
        WR_ADD(0) <= WRAD0_ipd;
    else
	WR_ADD <= x_add;
    end if;

   end process;

   wrapper_write_clk : process(WEN_ipd, WRCLK_ipd)

   begin
    if (WEN_ipd = '1') then
	WR_CLK <= WRCLK_ipd;
    else
	WR_CLK <= '0';
    end if;

   end process;

   process(WR_CLK)

    begin
      if WR_CLK = '1' then
        write_add(4) <= WRAD4_ipd;
        write_add(3) <= WRAD3_ipd;
        write_add(2) <= WRAD2_ipd;
        write_add(1) <= WRAD1_ipd;
        write_add(0) <= WRAD0_ipd;
      end if;

   end process;

   wrapper_write_data : process(WEN_ipd, WRDATA3_ipd, WRDATA2_ipd, WRDATA1_ipd, WRDATA0_ipd)

   begin
    if (WEN_ipd = '1') then
        DIN(3) <= WRDATA3_ipd;
        DIN(2) <= WRDATA2_ipd;
        DIN(1) <= WRDATA1_ipd;
        DIN(0) <= WRDATA0_ipd;
    else
	DIN <= x_data;
    end if;

   end process;


  VITALBehavior : PROCESS ( WEN_ipd, WR_CLK, DIN, RD_ADD, WR_ADD, WRAD4_ipd,WRAD3_ipd,WRAD2_ipd,WRAD1_ipd,WRAD0_ipd )


   -- Temporary variables
   VARIABLE tempaddr 		: integer := 0;
   VARIABLE rd_address 		: integer := 0;
   VARIABLE rd_viol_flag 	: X01 := '0';

   -- Timing Check results
   VARIABLE Pviol_WRCLK			: std_logic := '0';
   VARIABLE PeriodData_WRCLK		: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_WR_ADD_stp_hld_0	: std_logic := '0';
   VARIABLE TimingData_WR_ADD_stp_hld_0	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_WR_ADD_stp_hld_1	: std_logic := '0';
   VARIABLE TimingData_WR_ADD_stp_hld_1	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_WR_ADD_stp_hld_2	: std_logic := '0';
   VARIABLE TimingData_WR_ADD_stp_hld_2	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_WR_ADD_stp_hld_3	: std_logic := '0';
   VARIABLE TimingData_WR_ADD_stp_hld_3	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_WR_ADD_stp_hld_4	: std_logic := '0';
   VARIABLE TimingData_WR_ADD_stp_hld_4	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_WR_DATA_stp_0		: std_logic := '0';
   VARIABLE TimingData_WR_DATA_stp_0	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_WR_DATA_stp_1		: std_logic := '0';
   VARIABLE TimingData_WR_DATA_stp_1	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_WR_DATA_stp_2		: std_logic := '0';
   VARIABLE TimingData_WR_DATA_stp_2	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_WR_DATA_stp_3		: std_logic := '0';
   VARIABLE TimingData_WR_DATA_stp_3	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_WR_DATA_hld_0		: std_logic := '0';
   VARIABLE TimingData_WR_DATA_hld_0	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_WR_DATA_hld_1		: std_logic := '0';
   VARIABLE TimingData_WR_DATA_hld_1	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_WR_DATA_hld_2		: std_logic := '0';
   VARIABLE TimingData_WR_DATA_hld_2	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_WR_DATA_hld_3		: std_logic := '0';
   VARIABLE TimingData_WR_DATA_hld_3	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_WEN_stp_hld		: std_logic := '0';
   VARIABLE TimingData_WEN_stp_hld		: VitalTimingDataType := VitalTimingDataInit;



 BEGIN
    -------------------------------------------------------------------
    -- Timing Check Section
    -------------------------------------------------------------------
    IF (TimingChecksOn) THEN

	VitalPeriodPulseCheck  (Pviol_WRCLK,
				PeriodData_WRCLK,
				WR_CLK, "WRCLK",
				0.0 ns,
				0.0 ns,
				tpw_WRCLK_posedge,
				0.0 ns,
				TRUE,
				InstancePath & "/RB_MA",
				TRUE,
				TRUE,
				WARNING );

        VitalSetupHoldCheck    (Tviol_WR_ADD_stp_hld_0,
                                TimingData_WR_ADD_stp_hld_0,
                                WR_ADD(0), "WRAD0",
                                0.0 ns,
                                WR_CLK, "WRCLK",
                                0.0 ns,
                                tsetup_WRAD0_WRCLK_noedge_posedge, tsetup_WRAD0_WRCLK_noedge_posedge,
                                thold_WRAD0_WRCLK_noedge_posedge, thold_WRAD0_WRCLK_noedge_posedge,
                                WEN_ipd = '1',
                                '/',
                                InstancePath & "/RB_MA",
                                TRUE,
                                TRUE,
                                WARNING );

        VitalSetupHoldCheck    (Tviol_WR_ADD_stp_hld_1,
                                TimingData_WR_ADD_stp_hld_1,
                                WR_ADD(1), "WRAD1",
                                0.0 ns,
                                WR_CLK, "WRCLK",
                                0.0 ns,
                                tsetup_WRAD1_WRCLK_noedge_posedge, tsetup_WRAD1_WRCLK_noedge_posedge,
                                thold_WRAD1_WRCLK_noedge_posedge, thold_WRAD1_WRCLK_noedge_posedge,
                                WEN_ipd = '1',
                                '/',
                                InstancePath & "/RB_MA",
                                TRUE,
                                TRUE,
                                WARNING );

        VitalSetupHoldCheck    (Tviol_WR_ADD_stp_hld_2,
                                TimingData_WR_ADD_stp_hld_2,
                                WR_ADD(2), "WRAD2",
                                0.0 ns,
                                WR_CLK, "WRCLK",
                                0.0 ns,
                                tsetup_WRAD2_WRCLK_noedge_posedge, tsetup_WRAD2_WRCLK_noedge_posedge,
                                thold_WRAD2_WRCLK_noedge_posedge, thold_WRAD2_WRCLK_noedge_posedge,
                                WEN_ipd = '1',
                                '/',
                                InstancePath & "/RB_MA",
                                TRUE,
                                TRUE,
                                WARNING );

        VitalSetupHoldCheck    (Tviol_WR_ADD_stp_hld_3,
                                TimingData_WR_ADD_stp_hld_3,
                                WR_ADD(3), "WRAD3",
                                0.0 ns,
                                WR_CLK, "WRCLK",
                                0.0 ns,
                                tsetup_WRAD3_WRCLK_noedge_posedge, tsetup_WRAD3_WRCLK_noedge_posedge,
                                thold_WRAD3_WRCLK_noedge_posedge, thold_WRAD3_WRCLK_noedge_posedge,
                                WEN_ipd = '1',
                                '/',
                                InstancePath & "/RB_MA",
                                TRUE,
                                TRUE,
                                WARNING );
        VitalSetupHoldCheck    (Tviol_WR_ADD_stp_hld_4,
                                TimingData_WR_ADD_stp_hld_4,
                                WR_ADD(4), "WRAD4",
                                0.0 ns,
                                WR_CLK, "WRCLK",
                                0.0 ns,
                                tsetup_WRAD4_WRCLK_noedge_posedge, tsetup_WRAD4_WRCLK_noedge_posedge,
                                thold_WRAD4_WRCLK_noedge_posedge, thold_WRAD4_WRCLK_noedge_posedge,
                                WEN_ipd = '1',
                                '/',
                                InstancePath & "/RB_MA",
                                TRUE,
                                TRUE,
                                WARNING );

        VitalSetupHoldCheck    (Tviol_WR_DATA_stp_0,
                                TimingData_WR_DATA_stp_0,
                                DIN(0), "WRDATA0",
                                0.0 ns,
                                WR_CLK, "WRCLK",
                                0.0 ns,
                                tsetup_WRDATA0_WRCLK_noedge_posedge, tsetup_WRDATA0_WRCLK_noedge_posedge,
                                0.0 ns, 0.0 ns,
                                WEN_ipd = '1',
                                '/',
                                InstancePath & "/RB_MA",
                                TRUE,
                                TRUE,
                                WARNING );

        VitalSetupHoldCheck    (Tviol_WR_DATA_stp_1,
                                TimingData_WR_DATA_stp_1,
                                DIN(1), "WRDATA1",
                                0.0 ns,
                                WR_CLK, "WRCLK",
                                0.0 ns,
                                tsetup_WRDATA1_WRCLK_noedge_posedge, tsetup_WRDATA1_WRCLK_noedge_posedge,
                                0.0 ns, 0.0 ns,
                                WEN_ipd = '1',
                                '/',
                                InstancePath & "/RB_MA",
                                TRUE,
                                TRUE,
                                WARNING );

        VitalSetupHoldCheck    (Tviol_WR_DATA_stp_2,
                                TimingData_WR_DATA_stp_2,
                                DIN(2), "WRDATA2",
                                0.0 ns,
                                WR_CLK, "WRCLK",
                                0.0 ns,
                                tsetup_WRDATA2_WRCLK_noedge_posedge, tsetup_WRDATA2_WRCLK_noedge_posedge,
                                0.0 ns, 0.0 ns,
                                WEN_ipd = '1',
                                '/',
                                InstancePath & "/RB_MA",
                                TRUE,
                                TRUE,
                                WARNING );
        VitalSetupHoldCheck    (Tviol_WR_DATA_stp_3,
                                TimingData_WR_DATA_stp_3,
                                DIN(3), "WRDATA3",
                                0.0 ns,
                                WR_CLK, "WRCLK",
                                0.0 ns,
                                tsetup_WRDATA3_WRCLK_noedge_posedge, tsetup_WRDATA3_WRCLK_noedge_posedge,
                                0.0 ns, 0.0 ns,
                                WEN_ipd = '1',
                                '/',
                                InstancePath & "/RB_MA",
                                TRUE,
                                TRUE,
                                WARNING );

        VitalSetupHoldCheck    (Tviol_WR_DATA_hld_0,
                                TimingData_WR_DATA_hld_0,
                                DIN(0), "WRDATA0",
                                0.0 ns,
                                WR_CLK, "WRCLK",
                                0.0 ns,
                                0.0 ns, 0.0 ns,
                                thold_WRDATA0_WRCLK_noedge_posedge, thold_WRDATA0_WRCLK_noedge_posedge,
                                WEN_ipd = '1',
                                '/',
                                InstancePath & "/RB_MA",
                                TRUE,
                                TRUE,
                                WARNING );

        VitalSetupHoldCheck    (Tviol_WR_DATA_hld_1,
                                TimingData_WR_DATA_hld_1,
                                DIN(1), "WRDATA1",
                                0.0 ns,
                                WR_CLK, "WRCLK",
                                0.0 ns,
                                0.0 ns, 0.0 ns,
                                thold_WRDATA1_WRCLK_noedge_posedge, thold_WRDATA1_WRCLK_noedge_posedge,
                                WEN_ipd = '1',
                                '/',
                                InstancePath & "/RB_MA",
                                TRUE,
                                TRUE,
                                WARNING );

        VitalSetupHoldCheck    (Tviol_WR_DATA_hld_2,
                                TimingData_WR_DATA_hld_2,
                                DIN(2), "WRDATA2",
                                0.0 ns,
                                WR_CLK, "WRCLK",
                                0.0 ns,
                                0.0 ns, 0.0 ns,
                                thold_WRDATA2_WRCLK_noedge_posedge, thold_WRDATA2_WRCLK_noedge_posedge,
                                WEN_ipd = '1',
                                '/',
                                InstancePath & "/RB_MA",
                                TRUE,
                                TRUE,
                                WARNING );
        VitalSetupHoldCheck    (Tviol_WR_DATA_hld_3,
                                TimingData_WR_DATA_hld_3,
                                DIN(3), "WRDATA3",
                                0.0 ns,
                                WR_CLK, "WRCLK",
                                0.0 ns,
                                0.0 ns, 0.0 ns,
                                thold_WRDATA3_WRCLK_noedge_posedge, thold_WRDATA3_WRCLK_noedge_posedge,
                                WEN_ipd = '1',
                                '/',
                                InstancePath & "/RB_MA",
                                TRUE,
                                TRUE,
                                WARNING );


	VitalSetupHoldCheck    (Tviol_WEN_stp_hld,
				TimingData_WEN_stp_hld,
				WEN_ipd, "WEN",
				0.0 ns,
				WR_CLK, "WRCLK",
				0.0 ns,
				tsetup_WEN_WRCLK_noedge_posedge, tsetup_WEN_WRCLK_noedge_posedge,
				thold_WEN_WRCLK_noedge_posedge, thold_WEN_WRCLK_noedge_posedge,
				True,
				'/',
				InstancePath & "/RB_MA",
				TRUE,
				TRUE,
				WARNING );

    END IF; -- Timing Check Section


    -------------------------------------------------------------------
    -- Functionality Section
    -------------------------------------------------------------------

-- WRITE ADDRESS GOES XX

    if ( WR_CLK'EVENT and WR_CLK = '1' and vecX(WR_ADD)) then

        assert false
        report "Illegal Address Input: Undefined  Address at the Read_Write Port."
        severity note ;
        memory_array <= (others => x_data);

    end if;

-- ADDRESS HOLD AND SETUP VIOLATION EFFECT

    if( Tviol_WR_ADD_stp_hld_0 = 'X' or Tviol_WR_ADD_stp_hld_1 = 'X' or Tviol_WR_ADD_stp_hld_2 = 'X' or Tviol_WR_ADD_stp_hld_3 = 'X' or Tviol_WR_ADD_stp_hld_4 = 'X' ) then

        memory_array <= (others => x_data);

    else

-- DATA SETUP AND HOLD VIOLATION EFFECT

    if( Pviol_WRCLK = 'X' or Tviol_WR_DATA_hld_0 = 'X' or Tviol_WR_DATA_hld_1 = 'X' or Tviol_WR_DATA_hld_2 = 'X' or Tviol_WR_DATA_hld_3 = 'X' or Tviol_WEN_stp_hld = 'X') then
	tempaddr := vec2int(write_add);
	memory_array(tempaddr) <= x_data;
    end if;

    if( Tviol_WR_DATA_stp_0 = 'X' or Tviol_WR_DATA_stp_1 = 'X' or Tviol_WR_DATA_stp_2 = 'X' or Tviol_WR_DATA_stp_3 = 'X') then
	tempaddr := vec2int(WR_ADD);
	memory_array(tempaddr) <= x_data;
    end if;

    end if;

-- VALID MEMORY WRITE

    if ( WR_CLK'EVENT and WR_CLK = '1' and not(vecX(WR_ADD)) and not(Tviol_WR_ADD_stp_hld_0 = 'X' or Tviol_WR_ADD_stp_hld_1 = 'X' or Tviol_WR_ADD_stp_hld_2 = 'X' or Tviol_WR_ADD_stp_hld_3 = 'X' or Tviol_WR_ADD_stp_hld_4 = 'X') and not( Pviol_WRCLK = 'X' or Tviol_WR_DATA_hld_0 = 'X' or Tviol_WR_DATA_hld_1 = 'X' or Tviol_WR_DATA_hld_2 = 'X' or Tviol_WR_DATA_hld_3 = 'X' or Tviol_WEN_stp_hld = 'X') and not( Tviol_WR_DATA_stp_0 = 'X' or Tviol_WR_DATA_stp_1 = 'X' or Tviol_WR_DATA_stp_2 = 'X' or Tviol_WR_DATA_stp_3 = 'X')) then
	tempaddr := vec2int(WR_ADD);
	memory_array(tempaddr) <= DIN;
    end if;

    if WR_CLK'EVENT and WR_CLK /= WRCLK_ipd and WR_CLK'LAST_VALUE = '1' then
	memory_array(tempaddr) <= x_data;
    end if;


-- READ CYCLE VIOLATION EFFECT

    if(RD_ADD'EVENT and vecX(RD_ADD)) then
	data_out <= x_data;
    elsif

-- VALID MEMORY READ

     (RD_ADD'EVENT and not (vecX(RD_ADD))) then
	rd_address := vec2int(RD_ADD);
	data_out <= TRANSPORT memory_array(rd_address);
    end if;


  END PROCESS;

    -------------------------------------------------------------------------------
    -- Temporary output signal should get assigned to the output signal.
    -------------------------------------------------------------------------------

   PROCESS(data_out, OE_ipd, WRAD4_ipd,WRAD3_ipd,WRAD2_ipd,WRAD1_ipd,WRAD0_ipd)

   VARIABLE GLITCH_DATA : VitalGlitchDataType;
   VARIABLE con : std_logic := '0';
    VARIABLE WEN_inv : std_logic := '0';
    VARIABLE WRDATA3_1 : std_logic := 'Z';
    VARIABLE WRDATA2_1 : std_logic := 'Z';
    VARIABLE WRDATA1_1 : std_logic := 'Z';
    VARIABLE WRDATA0_1 : std_logic := 'Z';

   BEGIN
       WEN_inv := VitalINV(WEN_ipd);
       con := VitalAND2(OE_ipd,WEN_inv);


      WRDATA3_1 := VITALBUFIF1(data_out(3),con);
      WRDATA2_1 := VITALBUFIF1(data_out(2),con);
      WRDATA1_1 := VITALBUFIF1(data_out(1),con);
      WRDATA0_1 := VITALBUFIF1(data_out(0),con);

      VitalPathDelay01Z ( WRDATA3, GLITCH_DATA, "WRDATA3", WRDATA3_1,
        Paths => (
        0 => ( WRAD4_ipd'LAST_EVENT, VitalExtendToFillDelay(tpd_WRAD4_WRDATA3), TRUE ),
        1 => ( WRAD3_ipd'LAST_EVENT, VitalExtendToFillDelay(tpd_WRAD3_WRDATA3), TRUE ),
        2 => ( WRAD2_ipd'LAST_EVENT, VitalExtendToFillDelay(tpd_WRAD2_WRDATA3), TRUE ),
        3 => ( WRAD1_ipd'LAST_EVENT, VitalExtendToFillDelay(tpd_WRAD1_WRDATA3), TRUE ),
        4 => ( WRAD0_ipd'LAST_EVENT, VitalExtendToFillDelay(tpd_WRAD0_WRDATA3), TRUE ),
        5 => ( OE_ipd'LAST_EVENT, VitalExtendToFillDelay(tpd_OE_WRDATA3), TRUE ) ),
        DefaultDelay=>VitalZeroDelay01Z,
        Mode=>VitalInertial,
        XON=>TRUE,
        MsgOn=>TRUE,
        MsgSeverity=>WARNING,
        OutputMap => "UX01ZWLH-");

      VitalPathDelay01Z ( WRDATA2, GLITCH_DATA, "WRDATA2", WRDATA2_1,
        Paths => (
        0 => ( WRAD4_ipd'LAST_EVENT, VitalExtendToFillDelay(tpd_WRAD4_WRDATA2), TRUE ),
        1 => ( WRAD3_ipd'LAST_EVENT, VitalExtendToFillDelay(tpd_WRAD3_WRDATA2), TRUE ),
        2 => ( WRAD2_ipd'LAST_EVENT, VitalExtendToFillDelay(tpd_WRAD2_WRDATA2), TRUE ),
        3 => ( WRAD1_ipd'LAST_EVENT, VitalExtendToFillDelay(tpd_WRAD1_WRDATA2), TRUE ),
        4 => ( WRAD0_ipd'LAST_EVENT, VitalExtendToFillDelay(tpd_WRAD0_WRDATA2), TRUE ),
        5 => ( OE_ipd'LAST_EVENT, VitalExtendToFillDelay(tpd_OE_WRDATA2), TRUE ) ),
        DefaultDelay=>VitalZeroDelay01Z,
        Mode=>VitalInertial,
        XON=>TRUE,
        MsgOn=>TRUE,
        MsgSeverity=>WARNING,
        OutputMap => "UX01ZWLH-");

      VitalPathDelay01Z ( WRDATA1, GLITCH_DATA, "WRDATA1", WRDATA1_1,
        Paths => (
        0 => ( WRAD4_ipd'LAST_EVENT, VitalExtendToFillDelay(tpd_WRAD4_WRDATA1), TRUE ),
        1 => ( WRAD3_ipd'LAST_EVENT, VitalExtendToFillDelay(tpd_WRAD3_WRDATA1), TRUE ),
        2 => ( WRAD2_ipd'LAST_EVENT, VitalExtendToFillDelay(tpd_WRAD2_WRDATA1), TRUE ),
        3 => ( WRAD1_ipd'LAST_EVENT, VitalExtendToFillDelay(tpd_WRAD1_WRDATA1), TRUE ),
        4 => ( WRAD0_ipd'LAST_EVENT, VitalExtendToFillDelay(tpd_WRAD0_WRDATA1), TRUE ),
        5 => ( OE_ipd'LAST_EVENT, VitalExtendToFillDelay(tpd_OE_WRDATA1), TRUE ) ),
        DefaultDelay=>VitalZeroDelay01Z,
        Mode=>VitalInertial,
        XON=>TRUE,
        MsgOn=>TRUE,
        MsgSeverity=>WARNING,
        OutputMap => "UX01ZWLH-");

       VitalPathDelay01Z ( WRDATA0, GLITCH_DATA, "WRDATA0", WRDATA0_1,
        Paths => (
        0 => ( WRAD4_ipd'LAST_EVENT, VitalExtendToFillDelay(tpd_WRAD4_WRDATA0), TRUE ),
        1 => ( WRAD3_ipd'LAST_EVENT, VitalExtendToFillDelay(tpd_WRAD3_WRDATA0), TRUE ),
        2 => ( WRAD2_ipd'LAST_EVENT, VitalExtendToFillDelay(tpd_WRAD2_WRDATA0), TRUE ),
        3 => ( WRAD1_ipd'LAST_EVENT, VitalExtendToFillDelay(tpd_WRAD1_WRDATA0), TRUE ),
        4 => ( WRAD0_ipd'LAST_EVENT, VitalExtendToFillDelay(tpd_WRAD0_WRDATA0), TRUE ),
        5 => ( OE_ipd'LAST_EVENT, VitalExtendToFillDelay(tpd_OE_WRDATA0), TRUE ) ),
        DefaultDelay=>VitalZeroDelay01Z,
        Mode=>VitalInertial,
        XON=>TRUE,
        MsgOn=>TRUE,
        MsgSeverity=>WARNING,
        OutputMap => "UX01ZWLH-");

END PROCESS;

END VITAL_VF;
configuration CFG_RB_MA_VITAL of RB_MA is
        for VITAL_VF
        end for;
end CFG_RB_MA_VITAL;
-----------------------------------------------------------------------

-- VITAL model for RB_MS 30.10 technology
-----------------------------------------------------------------------

LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.VITAL_timing.all;
USE IEEE.VITAL_primitives.all;
LIBRARY VF1;
USE VF1.ALL;
USE VF1.RAMPACK.ALL;

-----------------------------------------------------------------------
-- ENTITY declaration
-----------------------------------------------------------------------

ENTITY RB_MS IS
  GENERIC (
	tipd_WEN		: VitalDelayType01			:= (0.0 ns, 0.0 ns);
	tipd_WRCLK		: VitalDelayType01			:= (0.0 ns, 0.0 ns);
	tipd_OE		: VitalDelayType01			:= (0.0 ns, 0.0 ns);
	tipd_WRDATA3		: VitalDelayType01	:= (0.0 ns, 0.0 ns);
	tipd_WRDATA2		: VitalDelayType01	:= (0.0 ns, 0.0 ns);
	tipd_WRDATA1		: VitalDelayType01	:= (0.0 ns, 0.0 ns);
	tipd_WRDATA0		: VitalDelayType01	:= (0.0 ns, 0.0 ns);
	tipd_WRAD4		: VitalDelayType01	:= (0.0 ns, 0.0 ns);
	tipd_WRAD3		: VitalDelayType01	:= (0.0 ns, 0.0 ns);
	tipd_WRAD2		: VitalDelayType01	:= (0.0 ns, 0.0 ns);
	tipd_WRAD1		: VitalDelayType01	:= (0.0 ns, 0.0 ns);
	tipd_WRAD0		: VitalDelayType01	:= (0.0 ns, 0.0 ns);

	tsetup_WRDATA3_WRCLK_noedge_posedge		: VitalDelayType :=  1 ns;
	tsetup_WRDATA2_WRCLK_noedge_posedge		: VitalDelayType :=  1 ns;
	tsetup_WRDATA1_WRCLK_noedge_posedge		: VitalDelayType :=  1 ns;
	tsetup_WRDATA0_WRCLK_noedge_posedge		: VitalDelayType :=  1 ns;
	tsetup_WRAD4_WRCLK_noedge_posedge		: VitalDelayType :=  1 ns;
	tsetup_WRAD3_WRCLK_noedge_posedge		: VitalDelayType :=  1 ns;
	tsetup_WRAD2_WRCLK_noedge_posedge		: VitalDelayType :=  1 ns;
	tsetup_WRAD1_WRCLK_noedge_posedge		: VitalDelayType :=  1 ns;
	tsetup_WRAD0_WRCLK_noedge_posedge		: VitalDelayType :=  1 ns;
	thold_WRDATA3_WRCLK_noedge_posedge		: VitalDelayType :=  1 ns;
	thold_WRDATA2_WRCLK_noedge_posedge		: VitalDelayType :=  1 ns;
	thold_WRDATA1_WRCLK_noedge_posedge		: VitalDelayType :=  1 ns;
	thold_WRDATA0_WRCLK_noedge_posedge		: VitalDelayType :=  1 ns;
	thold_WRAD4_WRCLK_noedge_posedge		: VitalDelayType :=  1 ns;
	thold_WRAD3_WRCLK_noedge_posedge		: VitalDelayType :=  1 ns;
	thold_WRAD2_WRCLK_noedge_posedge		: VitalDelayType :=  1 ns;
	thold_WRAD1_WRCLK_noedge_posedge		: VitalDelayType :=  1 ns;
	thold_WRAD0_WRCLK_noedge_posedge		: VitalDelayType :=  1 ns;
	tpw_WRCLK_posedge					: VitalDelayType := 1 ns;
	tsetup_WEN_WRCLK_noedge_posedge			: VitalDelayType := 1 ns;
	thold_WEN_WRCLK_noedge_posedge			: VitalDelayType := 1 ns;

	tpd_WRCLK_WRDATA3			: VitalDelayType01Z := (2 ns,2 ns,2 ns,2 ns,2 ns,2 ns);
	tpd_WRCLK_WRDATA2			: VitalDelayType01Z := (2 ns,2 ns,2 ns,2 ns,2 ns,2 ns);
	tpd_WRCLK_WRDATA1			: VitalDelayType01Z := (2 ns,2 ns,2 ns,2 ns,2 ns,2 ns);
	tpd_WRCLK_WRDATA0			: VitalDelayType01Z := (2 ns,2 ns,2 ns,2 ns,2 ns,2 ns);

	tpd_OE_WRDATA3			: VitalDelayType01Z := (2 ns,2 ns,2 ns,2 ns,2 ns,2 ns);
	tpd_OE_WRDATA2			: VitalDelayType01Z := (2 ns,2 ns,2 ns,2 ns,2 ns,2 ns);
	tpd_OE_WRDATA1			: VitalDelayType01Z := (2 ns,2 ns,2 ns,2 ns,2 ns,2 ns);
	tpd_OE_WRDATA0			: VitalDelayType01Z := (2 ns,2 ns,2 ns,2 ns,2 ns,2 ns);

	TimingChecksOn : BOOLEAN := TRUE;
	InstancePath : STRING := "*"
            );
  PORT	(
	WEN		: IN	std_logic ;
	WRCLK		: IN	std_logic ;
	OE		: IN	std_logic ;
	WRDATA3	: INOUT	std_logic := 'Z';
	WRDATA2	: INOUT	std_logic := 'Z';
	WRDATA1	: INOUT	std_logic := 'Z';
	WRDATA0	: INOUT	std_logic := 'Z';
	WRAD4		: IN	std_logic;
	WRAD3		: IN	std_logic;
	WRAD2		: IN	std_logic;
	WRAD1		: IN	std_logic;
	WRAD0		: IN	std_logic
	);


   ATTRIBUTE VITAL_LEVEL0 OF RB_MS : ENTITY IS TRUE;

END RB_MS;

-----------------------------------------------------------------------
-- ARCHITECTURE declaration
-----------------------------------------------------------------------
ARCHITECTURE VITAL_VF OF RB_MS IS

    ATTRIBUTE VITAL_LEVEL1 OF VITAL_VF : ARCHITECTURE IS FALSE;

	SIGNAL WEN_ipd		: std_logic := 'X';
	SIGNAL WRCLK_ipd		: std_logic := '0';
	SIGNAL WR_CLK		: std_logic := '0';
	SIGNAL RD_CLK		: std_logic := '0';
	SIGNAL OE_ipd	: std_logic := 'X';
	SIGNAL WRDATA3_ipd	: std_logic := 'Z';
	SIGNAL WRDATA2_ipd	: std_logic := 'Z';
	SIGNAL WRDATA1_ipd	: std_logic := 'Z';
	SIGNAL WRDATA0_ipd	: std_logic := 'Z';
	SIGNAL DIN		: std_logic_vector(3 DOWNTO 0);
	SIGNAL RD_ADD		: std_logic_vector(4 DOWNTO 0);
	SIGNAL WRAD4_ipd		: std_logic := '0';
	SIGNAL WRAD3_ipd		: std_logic := '0';
	SIGNAL WRAD2_ipd		: std_logic := '0';
	SIGNAL WRAD1_ipd		: std_logic := '0';
	SIGNAL WRAD0_ipd		: std_logic := '0';
	SIGNAL WR_ADD		: std_logic_vector(4 DOWNTO 0);
	SIGNAL write_add	: std_logic_vector(4 DOWNTO 0);
	SIGNAL data_out		: std_logic_vector(3 DOWNTO 0);
	SIGNAL output_delay	: time		:= 0 ns;

BEGIN
   
  ---------------------------------------------------------------------
  -- INPUT PATH DELAYs
  ---------------------------------------------------------------------
  WIREDELAY : BLOCK
  BEGIN
	VitalWireDelay (WEN_ipd,		WEN,		tipd_WEN);
	VitalWireDelay (WRCLK_ipd,		WRCLK,		tipd_WRCLK);
	VitalWireDelay (OE_ipd,		OE,		tipd_OE);
	VitalWireDelay (WRDATA0_ipd,	WRDATA0,	tipd_WRDATA0);
	VitalWireDelay (WRDATA1_ipd,	WRDATA1,	tipd_WRDATA1);
	VitalWireDelay (WRDATA2_ipd,	WRDATA2,	tipd_WRDATA2);
	VitalWireDelay (WRDATA3_ipd,	WRDATA3,	tipd_WRDATA3);
	VitalWireDelay (WRAD0_ipd,		WRAD0,		tipd_WRAD0);
	VitalWireDelay (WRAD1_ipd,		WRAD1,		tipd_WRAD1);
	VitalWireDelay (WRAD2_ipd,		WRAD2,		tipd_WRAD2);
	VitalWireDelay (WRAD3_ipd,		WRAD3,		tipd_WRAD3);
	VitalWireDelay (WRAD4_ipd,		WRAD4,		tipd_WRAD4);

  END BLOCK;

  ---------------------------------------------------------------------
  -- Behavior Section
  ---------------------------------------------------------------------

  ---------------------------------------------------------------------
  -- Wrapper Section
  ---------------------------------------------------------------------

   wrapper_read_add : process(OE_ipd, WRAD4_ipd,WRAD3_ipd,WRAD2_ipd,WRAD1_ipd,WRAD0_ipd, WEN_ipd)

   begin
    if (OE_ipd = '1' and WEN_ipd = '0') then
	RD_ADD(4) <= WRAD4_ipd;
	RD_ADD(3) <= WRAD3_ipd;
	RD_ADD(2) <= WRAD2_ipd;
	RD_ADD(1) <= WRAD1_ipd;
	RD_ADD(0) <= WRAD0_ipd;
    else
	RD_ADD <= x_add;
    end if;

   end process;

   wrapper_read_clk : process(OE_ipd, WRCLK_ipd, WEN_ipd)

   begin
    if (OE_ipd = '1' and WEN_ipd = '0') then
	RD_CLK <= WRCLK_ipd;
    else
	RD_CLK <= '0';
    end if;

   end process;

   wrapper_write_add : process(WEN_ipd, WRAD4_ipd,WRAD3_ipd,WRAD2_ipd,WRAD1_ipd,WRAD0_ipd)

   begin
    if (WEN_ipd = '1') then
	WR_ADD(4) <= WRAD4_ipd;
	WR_ADD(3) <= WRAD3_ipd;
	WR_ADD(2) <= WRAD2_ipd;
	WR_ADD(1) <= WRAD1_ipd;
	WR_ADD(0) <= WRAD0_ipd;
    else
	WR_ADD <= x_add;
    end if;

   end process;

   wrapper_write_clk : process(WEN_ipd, WRCLK_ipd)

   begin
    if (WEN_ipd = '1') then
	WR_CLK <= WRCLK_ipd;
    else
	WR_CLK <= '0';
    end if;

   end process;

   process(WR_CLK)

    begin
      if WR_CLK = '1' then
	write_add(4) <= WRAD4_ipd;
	write_add(3) <= WRAD3_ipd;
	write_add(2) <= WRAD2_ipd;
	write_add(1) <= WRAD1_ipd;
	write_add(0) <= WRAD0_ipd;
      end if;

   end process;

   wrapper_write_data : process(WEN_ipd, WRDATA3_ipd, WRDATA2_ipd, WRDATA1_ipd, WRDATA0_ipd)

   begin
    if (WEN_ipd = '1') then
	DIN(3) <= WRDATA3_ipd;
	DIN(2) <= WRDATA2_ipd;
	DIN(1) <= WRDATA1_ipd;
	DIN(0) <= WRDATA0_ipd;
    else
	DIN <= x_data;
    end if;

   end process;


  VITALBehavior : PROCESS ( WEN_ipd, write_add, WR_CLK, RD_CLK, DIN, RD_ADD, WR_ADD )

   VARIABLE memory_array : memory_array_typ;

   -- Temporary variables
   VARIABLE tempaddr : integer := 0;
   VARIABLE rd_address : integer := 0;

   -- Timing Check results
   VARIABLE Pviol_RDCLK			: std_logic := '0';
   VARIABLE PeriodData_RDCLK		: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_WRCLK			: std_logic := '0';
   VARIABLE PeriodData_WRCLK		: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_WR_ADD_stp_hld_0	: std_logic := '0';
   VARIABLE TimingData_WR_ADD_stp_hld_0	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_WR_ADD_stp_hld_1	: std_logic := '0';
   VARIABLE TimingData_WR_ADD_stp_hld_1	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_WR_ADD_stp_hld_2	: std_logic := '0';
   VARIABLE TimingData_WR_ADD_stp_hld_2	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_WR_ADD_stp_hld_3	: std_logic := '0';
   VARIABLE TimingData_WR_ADD_stp_hld_3	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_WR_ADD_stp_hld_4	: std_logic := '0';
   VARIABLE TimingData_WR_ADD_stp_hld_4	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_WR_DATA_stp_0		: std_logic := '0';
   VARIABLE TimingData_WR_DATA_stp_0	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_WR_DATA_stp_1		: std_logic := '0';
   VARIABLE TimingData_WR_DATA_stp_1	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_WR_DATA_stp_2		: std_logic := '0';
   VARIABLE TimingData_WR_DATA_stp_2	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_WR_DATA_stp_3		: std_logic := '0';
   VARIABLE TimingData_WR_DATA_stp_3	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_WR_DATA_hld_0		: std_logic := '0';
   VARIABLE TimingData_WR_DATA_hld_0	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_WR_DATA_hld_1		: std_logic := '0';
   VARIABLE TimingData_WR_DATA_hld_1	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_WR_DATA_hld_2		: std_logic := '0';
   VARIABLE TimingData_WR_DATA_hld_2	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_WR_DATA_hld_3		: std_logic := '0';
   VARIABLE TimingData_WR_DATA_hld_3	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_RD_ADD_stp_hld_0	: std_logic := '0';
   VARIABLE TimingData_RD_ADD_stp_hld_0	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_RD_ADD_stp_hld_1	: std_logic := '0';
   VARIABLE TimingData_RD_ADD_stp_hld_1	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_RD_ADD_stp_hld_2	: std_logic := '0';
   VARIABLE TimingData_RD_ADD_stp_hld_2	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_RD_ADD_stp_hld_3	: std_logic := '0';
   VARIABLE TimingData_RD_ADD_stp_hld_3	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_RD_ADD_stp_hld_4	: std_logic := '0';
   VARIABLE TimingData_RD_ADD_stp_hld_4	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_WEN_hld		: std_logic := '0';
   VARIABLE TimingData_WEN_hld		: VitalTimingDataType := VitalTimingDataInit;



 BEGIN
    -------------------------------------------------------------------
    -- Timing Check Section
    -------------------------------------------------------------------
    IF (TimingChecksOn) THEN

	VitalPeriodPulseCheck  (Pviol_RDCLK,
				PeriodData_RDCLK,
				RD_CLK, "WRCLK",
				0.0 ns,
				0.0 ns,
				tpw_WRCLK_posedge,
				0.0 ns,
				OE_ipd = '1' and WEN_ipd = '0',
				InstancePath & "/RB_MS",
				TRUE,
				TRUE,
				WARNING );

	VitalPeriodPulseCheck  (Pviol_WRCLK,
				PeriodData_WRCLK,
				WR_CLK, "WRCLK",
				0.0 ns,
				0.0 ns,
				tpw_WRCLK_posedge,
				0.0 ns,
				WEN_ipd = '1',
				InstancePath & "/RB_MS",
				TRUE,
				TRUE,
				WARNING );

	VitalSetupHoldCheck    (Tviol_WR_ADD_stp_hld_0,
				TimingData_WR_ADD_stp_hld_0,
				WR_ADD(0), "WRAD0",
				0.0 ns,
				WR_CLK, "WRCLK",
				0.0 ns,
				tsetup_WRAD0_WRCLK_noedge_posedge, tsetup_WRAD0_WRCLK_noedge_posedge, 
				thold_WRAD0_WRCLK_noedge_posedge, thold_WRAD0_WRCLK_noedge_posedge,
				WEN_ipd = '1',
				'/',
				InstancePath & "/RB_MS",
				TRUE,
				TRUE,
				WARNING );

	VitalSetupHoldCheck    (Tviol_WR_ADD_stp_hld_1,
				TimingData_WR_ADD_stp_hld_1,
				WR_ADD(1), "WRAD1",
				0.0 ns,
				WR_CLK, "WRCLK",
				0.0 ns,
				tsetup_WRAD1_WRCLK_noedge_posedge, tsetup_WRAD1_WRCLK_noedge_posedge, 
				thold_WRAD1_WRCLK_noedge_posedge, thold_WRAD1_WRCLK_noedge_posedge,
				WEN_ipd = '1',
				'/',
				InstancePath & "/RB_MS",
				TRUE,
				TRUE,
				WARNING );

	VitalSetupHoldCheck    (Tviol_WR_ADD_stp_hld_2,
				TimingData_WR_ADD_stp_hld_2,
				WR_ADD(2), "WRAD2",
				0.0 ns,
				WR_CLK, "WRCLK",
				0.0 ns,
				tsetup_WRAD2_WRCLK_noedge_posedge, tsetup_WRAD2_WRCLK_noedge_posedge, 
				thold_WRAD2_WRCLK_noedge_posedge, thold_WRAD2_WRCLK_noedge_posedge,
				WEN_ipd = '1',
				'/',
				InstancePath & "/RB_MS",
				TRUE,
				TRUE,
				WARNING );

	VitalSetupHoldCheck    (Tviol_WR_ADD_stp_hld_3,
				TimingData_WR_ADD_stp_hld_3,
				WR_ADD(3), "WRAD3",
				0.0 ns,
				WR_CLK, "WRCLK",
				0.0 ns,
				tsetup_WRAD3_WRCLK_noedge_posedge, tsetup_WRAD3_WRCLK_noedge_posedge, 
				thold_WRAD3_WRCLK_noedge_posedge, thold_WRAD3_WRCLK_noedge_posedge,
				WEN_ipd = '1',
				'/',
				InstancePath & "/RB_MS",
				TRUE,
				TRUE,
				WARNING );

	VitalSetupHoldCheck    (Tviol_WR_ADD_stp_hld_4,
				TimingData_WR_ADD_stp_hld_4,
				WR_ADD(4), "WRAD4",
				0.0 ns,
				WR_CLK, "WRCLK",
				0.0 ns,
				tsetup_WRAD4_WRCLK_noedge_posedge, tsetup_WRAD4_WRCLK_noedge_posedge, 
				thold_WRAD4_WRCLK_noedge_posedge, thold_WRAD4_WRCLK_noedge_posedge,
				WEN_ipd = '1',
				'/',
				InstancePath & "/RB_MS",
				TRUE,
				TRUE,
				WARNING );

	VitalSetupHoldCheck    (Tviol_WR_DATA_stp_0,
				TimingData_WR_DATA_stp_0,
				DIN(0), "WRDATA0",
				0.0 ns,
				WR_CLK, "WRCLK",
				0.0 ns,
				tsetup_WRDATA0_WRCLK_noedge_posedge, tsetup_WRDATA0_WRCLK_noedge_posedge, 
				0.0 ns, 0.0 ns,
				WEN_ipd = '1',
				'/',
				InstancePath & "/RB_MS",
				TRUE,
				TRUE,
				WARNING );

	VitalSetupHoldCheck    (Tviol_WR_DATA_stp_1,
				TimingData_WR_DATA_stp_1,
				DIN(1), "WRDATA1",
				0.0 ns,
				WR_CLK, "WRCLK",
				0.0 ns,
				tsetup_WRDATA1_WRCLK_noedge_posedge, tsetup_WRDATA1_WRCLK_noedge_posedge, 
				0.0 ns, 0.0 ns,
				WEN_ipd = '1',
				'/',
				InstancePath & "/RB_MS",
				TRUE,
				TRUE,
				WARNING );

	VitalSetupHoldCheck    (Tviol_WR_DATA_stp_2,
				TimingData_WR_DATA_stp_2,
				DIN(2), "WRDATA2",
				0.0 ns,
				WR_CLK, "WRCLK",
				0.0 ns,
				tsetup_WRDATA2_WRCLK_noedge_posedge, tsetup_WRDATA2_WRCLK_noedge_posedge, 
				0.0 ns, 0.0 ns,
				WEN_ipd = '1',
				'/',
				InstancePath & "/RB_MS",
				TRUE,
				TRUE,
				WARNING );

	VitalSetupHoldCheck    (Tviol_WR_DATA_stp_3,
				TimingData_WR_DATA_stp_3,
				DIN(3), "WRDATA3",
				0.0 ns,
				WR_CLK, "WRCLK",
				0.0 ns,
				tsetup_WRDATA3_WRCLK_noedge_posedge, tsetup_WRDATA3_WRCLK_noedge_posedge, 
				0.0 ns, 0.0 ns,
				WEN_ipd = '1',
				'/',
				InstancePath & "/RB_MS",
				TRUE,
				TRUE,
				WARNING );

	VitalSetupHoldCheck    (Tviol_WR_DATA_hld_0,
				TimingData_WR_DATA_hld_0,
				DIN(0), "WRDATA0",
				0.0 ns,
				WR_CLK, "WRCLK",
				0.0 ns,
				0.0 ns, 0.0 ns,
				thold_WRDATA0_WRCLK_noedge_posedge, thold_WRDATA0_WRCLK_noedge_posedge,
				WEN_ipd = '1',
				'/',
				InstancePath & "/RB_MS",
				TRUE,
				TRUE,
				WARNING );

	VitalSetupHoldCheck    (Tviol_WR_DATA_hld_1,
				TimingData_WR_DATA_hld_1,
				DIN(1), "WRDATA1",
				0.0 ns,
				WR_CLK, "WRCLK",
				0.0 ns,
				0.0 ns, 0.0 ns,
				thold_WRDATA1_WRCLK_noedge_posedge, thold_WRDATA1_WRCLK_noedge_posedge,
				WEN_ipd = '1',
				'/',
				InstancePath & "/RB_MS",
				TRUE,
				TRUE,
				WARNING );

	VitalSetupHoldCheck    (Tviol_WR_DATA_hld_2,
				TimingData_WR_DATA_hld_2,
				DIN(2), "WRDATA2",
				0.0 ns,
				WR_CLK, "WRCLK",
				0.0 ns,
				0.0 ns, 0.0 ns,
				thold_WRDATA2_WRCLK_noedge_posedge, thold_WRDATA2_WRCLK_noedge_posedge,
				WEN_ipd = '1',
				'/',
				InstancePath & "/RB_MS",
				TRUE,
				TRUE,
				WARNING );

	VitalSetupHoldCheck    (Tviol_WR_DATA_hld_3,
				TimingData_WR_DATA_hld_3,
				DIN(3), "WRDATA3",
				0.0 ns,
				WR_CLK, "WRCLK",
				0.0 ns,
				0.0 ns, 0.0 ns,
				thold_WRDATA3_WRCLK_noedge_posedge, thold_WRDATA3_WRCLK_noedge_posedge,
				WEN_ipd = '1',
				'/',
				InstancePath & "/RB_MS",
				TRUE,
				TRUE,
				WARNING );

	VitalSetupHoldCheck    (Tviol_RD_ADD_stp_hld_0,
				TimingData_RD_ADD_stp_hld_0,
				RD_ADD(0), "WRAD0",
				0.0 ns,
				RD_CLK, "WRCLK",
				0.0 ns,
				tsetup_WRAD0_WRCLK_noedge_posedge, tsetup_WRAD0_WRCLK_noedge_posedge, 
				thold_WRAD0_WRCLK_noedge_posedge, thold_WRAD0_WRCLK_noedge_posedge,
				OE_ipd = '1' and WEN_ipd = '0',
				'/',
				InstancePath & "/RB_MS",
				TRUE,
				TRUE,
				WARNING );

	VitalSetupHoldCheck    (Tviol_RD_ADD_stp_hld_1,
				TimingData_RD_ADD_stp_hld_1,
				RD_ADD(1), "WRAD1",
				0.0 ns,
				RD_CLK, "WRCLK",
				0.0 ns,
				tsetup_WRAD1_WRCLK_noedge_posedge, tsetup_WRAD1_WRCLK_noedge_posedge, 
				thold_WRAD1_WRCLK_noedge_posedge, thold_WRAD1_WRCLK_noedge_posedge,
				OE_ipd = '1' and WEN_ipd = '0',
				'/',
				InstancePath & "/RB_MS",
				TRUE,
				TRUE,
				WARNING );

	VitalSetupHoldCheck    (Tviol_RD_ADD_stp_hld_2,
				TimingData_RD_ADD_stp_hld_2,
				RD_ADD(2), "WRAD2",
				0.0 ns,
				RD_CLK, "WRCLK",
				0.0 ns,
				tsetup_WRAD2_WRCLK_noedge_posedge, tsetup_WRAD2_WRCLK_noedge_posedge, 
				thold_WRAD2_WRCLK_noedge_posedge, thold_WRAD2_WRCLK_noedge_posedge,
				OE_ipd = '1' and WEN_ipd = '0',
				'/',
				InstancePath & "/RB_MS",
				TRUE,
				TRUE,
				WARNING );

	VitalSetupHoldCheck    (Tviol_RD_ADD_stp_hld_3,
				TimingData_RD_ADD_stp_hld_3,
				RD_ADD(3), "WRAD3",
				0.0 ns,
				RD_CLK, "WRCLK",
				0.0 ns,
				tsetup_WRAD3_WRCLK_noedge_posedge, tsetup_WRAD3_WRCLK_noedge_posedge, 
				thold_WRAD3_WRCLK_noedge_posedge, thold_WRAD3_WRCLK_noedge_posedge,
				OE_ipd = '1' and WEN_ipd = '0',
				'/',
				InstancePath & "/RB_MS",
				TRUE,
				TRUE,
				WARNING );

	VitalSetupHoldCheck    (Tviol_RD_ADD_stp_hld_4,
				TimingData_RD_ADD_stp_hld_4,
				RD_ADD(4), "WRAD4",
				0.0 ns,
				RD_CLK, "WRCLK",
				0.0 ns,
				tsetup_WRAD4_WRCLK_noedge_posedge, tsetup_WRAD4_WRCLK_noedge_posedge, 
				thold_WRAD4_WRCLK_noedge_posedge, thold_WRAD4_WRCLK_noedge_posedge,
				OE_ipd = '1' and WEN_ipd = '0',
				'/',
				InstancePath & "/RB_MS",
				TRUE,
				TRUE,
				WARNING );

	VitalSetupHoldCheck    (Tviol_WEN_hld,
				TimingData_WEN_hld,
				WEN_ipd, "WEN",
				0.0 ns,
				WR_CLK, "WRCLK",
				0.0 ns,
				tsetup_WEN_WRCLK_noedge_posedge,tsetup_WEN_WRCLK_noedge_posedge,
				thold_WEN_WRCLK_noedge_posedge, thold_WEN_WRCLK_noedge_posedge,
				True,
				'/',
				InstancePath & "/RB_MS",
				TRUE,
				TRUE,
				WARNING );

    END IF; -- Timing Check Section

    -------------------------------------------------------------------
    -- Functionality Section
    -------------------------------------------------------------------

-- WRITE ADDRESS GOES XX

    if ( WR_CLK'EVENT and WR_CLK = '1' and vecX(WR_ADD)) then

        assert false
        report "Illegal Address Input: Undefined  Address at the Read_Write Port."
        severity note ;
        memory_array := (others => x_data);

    end if;

-- ADDRESS HOLD AND SETUP VIOLATION EFFECT

    if( Tviol_WR_ADD_stp_hld_0 = 'X' or Tviol_WR_ADD_stp_hld_1 = 'X' or Tviol_WR_ADD_stp_hld_2 = 'X' or Tviol_WR_ADD_stp_hld_3 = 'X' or Tviol_WR_ADD_stp_hld_4 = 'X' ) then
	memory_array := (others => x_data);
    else

-- DATA SETUP AND HOLD VIOLATION EFFECT

    if( Pviol_WRCLK = 'X' or Tviol_WR_DATA_hld_0 = 'X' or Tviol_WR_DATA_hld_1 = 'X' or Tviol_WR_DATA_hld_2 = 'X' or Tviol_WR_DATA_hld_3 = 'X' or Tviol_WEN_hld = 'X') then
	tempaddr := vec2int(write_add);
	memory_array(tempaddr) := x_data;
    end if;

    if( Tviol_WR_DATA_stp_0 = 'X' or Tviol_WR_DATA_stp_1 = 'X' or Tviol_WR_DATA_stp_2 = 'X' or Tviol_WR_DATA_stp_3 = 'X') then
	tempaddr := vec2int(write_add);
	memory_array(tempaddr) := x_data;
    end if;

    end if;

-- VALID MEMORY WRITE

    if ( WR_CLK'EVENT and WR_CLK = '1' and not(vecX(WR_ADD)) and not(Tviol_WR_ADD_stp_hld_0 = 'X' or Tviol_WR_ADD_stp_hld_1 = 'X' or Tviol_WR_ADD_stp_hld_2 = 'X' or Tviol_WR_ADD_stp_hld_3 = 'X' or Tviol_WR_ADD_stp_hld_4 = 'X' ) and not ( Pviol_WRCLK = 'X' or Tviol_WR_DATA_hld_0 = 'X' or Tviol_WR_DATA_hld_1 = 'X' or Tviol_WR_DATA_hld_2 = 'X' or Tviol_WR_DATA_hld_3 = 'X' or Tviol_WEN_hld = 'X') and not( Tviol_WR_DATA_stp_0 = 'X' or Tviol_WR_DATA_stp_1 = 'X' or Tviol_WR_DATA_stp_2 = 'X' or Tviol_WR_DATA_stp_3 = 'X')) then
	tempaddr := vec2int(WR_ADD);
	memory_array(tempaddr) := DIN;
    end if;

    if WR_CLK'EVENT and WR_CLK /= WRCLK_ipd and WR_CLK'LAST_VALUE = '1' then
	memory_array(tempaddr) := x_data;
    end if;


-- READ ADDRESS CYCLE VIOLATION EFFECT

    if( Tviol_RD_ADD_stp_hld_0 = 'X' or Tviol_RD_ADD_stp_hld_1 = 'X' or Tviol_RD_ADD_stp_hld_2 = 'X' or Tviol_RD_ADD_stp_hld_3 = 'X' or Tviol_RD_ADD_stp_hld_4 = 'X' or Pviol_RDCLK = 'X' or (RD_CLK'EVENT and RD_CLK = '1' and vecX(RD_ADD))) then
	--output_delay <= 0 ns;
	data_out <= x_data;
    elsif

-- VALID MEMORY READ

    (RD_CLK'EVENT and RD_CLK = '1' and not( Tviol_RD_ADD_stp_hld_0 = 'X' or Tviol_RD_ADD_stp_hld_1 = 'X' or Tviol_RD_ADD_stp_hld_2 = 'X' or Tviol_RD_ADD_stp_hld_3 = 'X' or Tviol_RD_ADD_stp_hld_4 = 'X' or Pviol_RDCLK = 'X' or vecX(RD_ADD) ))then
	rd_address := vec2int(RD_ADD);
	data_out <= memory_array(rd_address);
    end if;

    if RD_CLK'EVENT and RD_CLK /= WRCLK_ipd and RD_CLK'LAST_VALUE = '1' then
	--output_delay <= 0 ns;
	data_out <= x_data;
    end if;
     --data_out <= NULL;


  END PROCESS;

    -------------------------------------------------------------------------------
    -- Temporary output signal should get assigned to the output signal.
    -------------------------------------------------------------------------------

  PROCESS(data_out, WRCLK_ipd, WEN_ipd, OE_ipd)

    VARIABLE con : std_logic := '0';
    VARIABLE WEN_inv : std_logic := '0';
    VARIABLE WRDATA3_1 : std_logic := 'Z';
    VARIABLE WRDATA2_1 : std_logic := 'Z';
    VARIABLE WRDATA1_1 : std_logic := 'Z';
    VARIABLE WRDATA0_1 : std_logic := 'Z';
    VARIABLE GLITCH_DATA : VitalGlitchDataType;
    --VARIABLE GLITCH_DATA1 : VitalGlitchDataType;
    BEGIN
       
      WEN_inv := VitalINV(WEN_ipd);
      con := VitalAND2(WEN_inv,OE_ipd);
      WRDATA3_1 := VITALBUFIF1(data_out(3),con);
      WRDATA2_1 := VITALBUFIF1(data_out(2),con);
      WRDATA1_1 := VITALBUFIF1(data_out(1),con);
      WRDATA0_1 := VITALBUFIF1(data_out(0),con);

     VitalPathDelay01Z ( WRDATA3, GLITCH_DATA, "WRDATA3", WRDATA3_1,
        Paths => (
        0 => ( WRCLK_ipd'LAST_EVENT, VitalExtendToFillDelay(tpd_WRCLK_WRDATA3), TRUE ),
        1 => ( OE_ipd'LAST_EVENT, VitalExtendToFillDelay(tpd_OE_WRDATA3), TRUE ) ),
        DefaultDelay=>VitalZeroDelay01Z,
        Mode=>VitalInertial,
        XON=>TRUE,
        MsgOn=>TRUE,
        MsgSeverity=>WARNING, 
        OutputMap => "UX01ZWLH-");

     VitalPathDelay01Z ( WRDATA2, GLITCH_DATA, "WRDATA2", WRDATA2_1,
        Paths => (
        0 => ( WRCLK_ipd'LAST_EVENT, VitalExtendToFillDelay(tpd_WRCLK_WRDATA2), TRUE ),
        1 => ( OE_ipd'LAST_EVENT, VitalExtendToFillDelay(tpd_OE_WRDATA2), TRUE ) ),
        DefaultDelay=>VitalZeroDelay01Z,
        Mode=>VitalInertial,
        XON=>TRUE,
        MsgOn=>TRUE,
        MsgSeverity=>WARNING, 
        OutputMap => "UX01ZWLH-");

     VitalPathDelay01Z ( WRDATA1, GLITCH_DATA, "WRDATA1", WRDATA1_1,
        Paths => (
        0 => ( WRCLK_ipd'LAST_EVENT, VitalExtendToFillDelay(tpd_WRCLK_WRDATA1), TRUE ),
        1 => ( OE_ipd'LAST_EVENT, VitalExtendToFillDelay(tpd_OE_WRDATA1), TRUE ) ),
        DefaultDelay=>VitalZeroDelay01Z,
        Mode=>VitalInertial,
        XON=>TRUE,
        MsgOn=>TRUE,
        MsgSeverity=>WARNING, 
        OutputMap => "UX01ZWLH-");

     VitalPathDelay01Z ( WRDATA0, GLITCH_DATA, "WRDATA0", WRDATA0_1,
        Paths => (
        0 => ( WRCLK_ipd'LAST_EVENT, VitalExtendToFillDelay(tpd_WRCLK_WRDATA0), TRUE ),
        1 => ( OE_ipd'LAST_EVENT, VitalExtendToFillDelay(tpd_OE_WRDATA0), TRUE ))  ,
        DefaultDelay=>VitalZeroDelay01Z,
        Mode=>VitalInertial,
        XON=>TRUE,
        MsgOn=>TRUE,
        MsgSeverity=>WARNING, 
        OutputMap => "UX01ZWLH-");

END PROCESS;
END VITAL_VF;
configuration CFG_RB_MS_VITAL of RB_MS is
        for VITAL_VF
        end for;
end CFG_RB_MS_VITAL;
-----------------------------------------------------------------------

-- VITAL model for RB_SA 30.10 technology
-----------------------------------------------------------------------

LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.VITAL_timing.all;
USE IEEE.VITAL_primitives.all;
LIBRARY VF1;
USE VF1.ALL;
USE VF1.RAMPACK.ALL;

-----------------------------------------------------------------------
-- ENTITY declaration
-----------------------------------------------------------------------

ENTITY RB_SA IS
  GENERIC (
	tipd_WEN		: VitalDelayType01			:= (0.0 ns, 0.0 ns);
	tipd_REN		: VitalDelayType01			:= (0.0 ns, 0.0 ns);
	tipd_WCLK		: VitalDelayType01			:= (0.0 ns, 0.0 ns);
	tipd_WDATA3		: VitalDelayType01	                := (0.0 ns, 0.0 ns);
	tipd_WDATA2		: VitalDelayType01	                := (0.0 ns, 0.0 ns);
	tipd_WDATA1		: VitalDelayType01	                := (0.0 ns, 0.0 ns);
	tipd_WDATA0		: VitalDelayType01	                := (0.0 ns, 0.0 ns);
	tipd_RAD4		: VitalDelayType01	                := (0.0 ns, 0.0 ns);
	tipd_RAD3		: VitalDelayType01	                := (0.0 ns, 0.0 ns);
	tipd_RAD2		: VitalDelayType01	                := (0.0 ns, 0.0 ns);
	tipd_RAD1		: VitalDelayType01	                := (0.0 ns, 0.0 ns);
	tipd_RAD0		: VitalDelayType01	                := (0.0 ns, 0.0 ns);
	tipd_WAD4		: VitalDelayType01	                := (0.0 ns, 0.0 ns);
	tipd_WAD3		: VitalDelayType01	                := (0.0 ns, 0.0 ns);
	tipd_WAD2		: VitalDelayType01	                := (0.0 ns, 0.0 ns);
	tipd_WAD1		: VitalDelayType01	                := (0.0 ns, 0.0 ns);
	tipd_WAD0		: VitalDelayType01	                := (0.0 ns, 0.0 ns);

	tsetup_WDATA3_WCLK_noedge_posedge		: VitalDelayType := 1 ns;
	tsetup_WDATA2_WCLK_noedge_posedge		: VitalDelayType := 1 ns;
	tsetup_WDATA1_WCLK_noedge_posedge		: VitalDelayType := 1 ns;
	tsetup_WDATA0_WCLK_noedge_posedge		: VitalDelayType := 1 ns;

	thold_WDATA3_WCLK_noedge_posedge		: VitalDelayType := 1 ns;
	thold_WDATA2_WCLK_noedge_posedge		: VitalDelayType := 1 ns;
	thold_WDATA1_WCLK_noedge_posedge		: VitalDelayType := 1 ns;
	thold_WDATA0_WCLK_noedge_posedge		: VitalDelayType := 1 ns;

	tsetup_WAD4_WCLK_noedge_posedge		: VitalDelayType := 1 ns;
	tsetup_WAD3_WCLK_noedge_posedge		: VitalDelayType := 1 ns;
	tsetup_WAD2_WCLK_noedge_posedge		: VitalDelayType := 1 ns;
	tsetup_WAD1_WCLK_noedge_posedge		: VitalDelayType := 1 ns;
	tsetup_WAD0_WCLK_noedge_posedge		: VitalDelayType := 1 ns;

	thold_WAD4_WCLK_noedge_posedge		: VitalDelayType := 1 ns;
	thold_WAD3_WCLK_noedge_posedge		: VitalDelayType := 1 ns;
	thold_WAD2_WCLK_noedge_posedge		: VitalDelayType := 1 ns;
	thold_WAD1_WCLK_noedge_posedge		: VitalDelayType := 1 ns;
	thold_WAD0_WCLK_noedge_posedge		: VitalDelayType := 1 ns;

	tpw_WCLK_posedge              			: VitalDelayType			:= 1 ns;
	tsetup_WEN_WCLK_noedge_posedge		: VitalDelayType 			:= 1 ns;
	thold_WEN_WCLK_noedge_posedge		: VitalDelayType 			:= 1 ns;

        tpd_RAD4_RDATA0         :VitalDelayType01 := (2.0 ns,2.0 ns);
        tpd_RAD3_RDATA0         :VitalDelayType01 := (2.0 ns,2.0 ns);
        tpd_RAD2_RDATA0         :VitalDelayType01 := (2.0 ns,2.0 ns);
        tpd_RAD1_RDATA0         :VitalDelayType01 := (2.0 ns,2.0 ns);
        tpd_RAD0_RDATA0         :VitalDelayType01 := (2.0 ns,2.0 ns);
        tpd_RAD4_RDATA1         :VitalDelayType01 := (2.0 ns,2.0 ns);
        tpd_RAD3_RDATA1         :VitalDelayType01 := (2.0 ns,2.0 ns);
        tpd_RAD2_RDATA1         :VitalDelayType01 := (2.0 ns,2.0 ns);
        tpd_RAD1_RDATA1         :VitalDelayType01 := (2.0 ns,2.0 ns);
        tpd_RAD0_RDATA1         :VitalDelayType01 := (2.0 ns,2.0 ns);
        tpd_RAD4_RDATA2         :VitalDelayType01 := (2.0 ns,2.0 ns);
        tpd_RAD3_RDATA2         :VitalDelayType01 := (2.0 ns,2.0 ns);
        tpd_RAD2_RDATA2         :VitalDelayType01 := (2.0 ns,2.0 ns);
        tpd_RAD1_RDATA2         :VitalDelayType01 := (2.0 ns,2.0 ns);
        tpd_RAD0_RDATA2         :VitalDelayType01 := (2.0 ns,2.0 ns);
        tpd_RAD4_RDATA3         :VitalDelayType01 := (2.0 ns,2.0 ns);
        tpd_RAD3_RDATA3         :VitalDelayType01 := (2.0 ns,2.0 ns);
        tpd_RAD2_RDATA3         :VitalDelayType01 := (2.0 ns,2.0 ns);
        tpd_RAD1_RDATA3         :VitalDelayType01 := (2.0 ns,2.0 ns);
        tpd_RAD0_RDATA3         :VitalDelayType01 := (2.0 ns,2.0 ns);
        tpd_REN_RDATA0         :VitalDelayType01 := (2.0 ns,2.0 ns);
        tpd_REN_RDATA1         :VitalDelayType01 := (2.0 ns,2.0 ns);
        tpd_REN_RDATA2         :VitalDelayType01 := (2.0 ns,2.0 ns);
        tpd_REN_RDATA3         :VitalDelayType01 := (2.0 ns,2.0 ns);

	TimingChecksOn : BOOLEAN := TRUE;
	InstancePath : STRING := "*"
            );
  PORT	(
	WEN		: IN	std_logic ;
	REN		: IN	std_logic ;
	WCLK		: IN	std_logic ;
	WDATA3	        : IN	std_logic ;
	WDATA2	        : IN	std_logic ;
	WDATA1	        : IN	std_logic ;
	WDATA0	        : IN	std_logic ;
	RDATA3	        : OUT	std_logic ;
	RDATA2	        : OUT	std_logic ;
	RDATA1	        : OUT	std_logic ;
	RDATA0	        : OUT	std_logic ;
	RAD4		: IN	std_logic ;
	RAD3		: IN	std_logic ;
	RAD2		: IN	std_logic ;
	RAD1		: IN	std_logic ;
	RAD0		: IN	std_logic ;
	WAD4		: IN	std_logic ;
	WAD3		: IN	std_logic ;
	WAD2		: IN	std_logic ;
	WAD1		: IN	std_logic ;
	WAD0		: IN	std_logic 
	);


   ATTRIBUTE VITAL_LEVEL0 OF RB_SA : ENTITY IS TRUE;

END RB_SA;

-----------------------------------------------------------------------
-- ARCHITECTURE declaration
-----------------------------------------------------------------------
ARCHITECTURE VITAL_VF OF RB_SA IS

    ATTRIBUTE VITAL_LEVEL1 OF VITAL_VF : ARCHITECTURE IS FALSE;

	SIGNAL WEN_ipd		: std_logic := 'X';
	SIGNAL REN_ipd		: std_logic := 'X';
	SIGNAL WCLK_ipd		: std_logic := '0';
	SIGNAL WR_CLK		: std_logic := '0';
	SIGNAL WDATA3_ipd	: std_logic := 'Z';
	SIGNAL WDATA2_ipd	: std_logic := 'Z';
	SIGNAL WDATA1_ipd	: std_logic := 'Z';
	SIGNAL WDATA0_ipd	: std_logic := 'Z';
	SIGNAL DIN		: std_logic_vector(3 DOWNTO 0);
	SIGNAL RAD4_ipd		: std_logic ;
	SIGNAL RAD3_ipd		: std_logic ;
	SIGNAL RAD2_ipd		: std_logic ;
	SIGNAL RAD1_ipd		: std_logic ;
	SIGNAL RAD0_ipd		: std_logic ;
	SIGNAL RD_ADD		: std_logic_vector(4 DOWNTO 0);
	SIGNAL WAD4_ipd		: std_logic ;
	SIGNAL WAD3_ipd		: std_logic ;
	SIGNAL WAD2_ipd		: std_logic ;
	SIGNAL WAD1_ipd		: std_logic ;
	SIGNAL WAD0_ipd		: std_logic ;
	SIGNAL WR_ADD		: std_logic_vector(4 DOWNTO 0);
	SIGNAL write_add	: std_logic_vector(4 DOWNTO 0);
	SIGNAL data_out		: std_logic_vector(3 DOWNTO 0) := x_data;
        SIGNAL memory_array : memory_array_typ := (others => x_data);

BEGIN
   
  ---------------------------------------------------------------------
  -- INPUT PATH DELAYs
  ---------------------------------------------------------------------
  WIREDELAY : BLOCK
  BEGIN
	VitalWireDelay (WEN_ipd,		WEN,		tipd_WEN);
	VitalWireDelay (REN_ipd,		REN,		tipd_REN);
	VitalWireDelay (WCLK_ipd,		WCLK,		tipd_WCLK);
	VitalWireDelay (WDATA0_ipd,	        WDATA0,	        tipd_WDATA0);
	VitalWireDelay (WDATA1_ipd,	        WDATA1,	        tipd_WDATA1);
	VitalWireDelay (WDATA2_ipd,	        WDATA2,	        tipd_WDATA2);
	VitalWireDelay (WDATA3_ipd,	        WDATA3,	        tipd_WDATA3);
	VitalWireDelay (RAD0_ipd,		RAD0,		tipd_RAD0);
	VitalWireDelay (RAD1_ipd,		RAD1,		tipd_RAD1);
	VitalWireDelay (RAD2_ipd,		RAD2,		tipd_RAD2);
	VitalWireDelay (RAD3_ipd,		RAD3,		tipd_RAD3);
	VitalWireDelay (RAD4_ipd,		RAD4,		tipd_RAD4);
	VitalWireDelay (WAD0_ipd,		WAD0,		tipd_WAD0);
	VitalWireDelay (WAD1_ipd,		WAD1,		tipd_WAD1);
	VitalWireDelay (WAD2_ipd,		WAD2,		tipd_WAD2);
	VitalWireDelay (WAD3_ipd,		WAD3,		tipd_WAD3);
	VitalWireDelay (WAD4_ipd,		WAD4,		tipd_WAD4);

  END BLOCK;

  ---------------------------------------------------------------------
  -- Behavior Section
  ---------------------------------------------------------------------

  ---------------------------------------------------------------------
  -- Wrapper Section
  ---------------------------------------------------------------------

   wrapper_read_add : process(REN_ipd, RAD4_ipd, RAD3_ipd, RAD2_ipd, RAD1_ipd, RAD0_ipd)

   begin
    if (REN_ipd = '1') then
	RD_ADD(4) <= RAD4_ipd;
	RD_ADD(3) <= RAD3_ipd;
	RD_ADD(2) <= RAD2_ipd;
	RD_ADD(1) <= RAD1_ipd;
	RD_ADD(0) <= RAD0_ipd;
    else
	RD_ADD <= x_add;
    end if;

   end process;


   wrapper_write_add : process(WEN_ipd, WAD4_ipd, WAD3_ipd, WAD2_ipd, WAD1_ipd, WAD0_ipd)

   begin
    if (WEN_ipd = '1') then
	WR_ADD(4) <= WAD4_ipd;
	WR_ADD(3) <= WAD3_ipd;
	WR_ADD(2) <= WAD2_ipd;
	WR_ADD(1) <= WAD1_ipd;
	WR_ADD(0) <= WAD0_ipd;
    else
	WR_ADD <= x_add;
    end if;

   end process;

   wrapper_write_clk : process(WEN_ipd, WCLK_ipd)

   begin
    if (WEN_ipd = '1') then
	WR_CLK <= WCLK_ipd;
    else
	WR_CLK <= '0';
    end if;

   end process;

   process(WR_CLK)

    begin
      if WR_CLK = '1' then
	write_add(4) <= WAD4_ipd;
	write_add(3) <= WAD3_ipd;
	write_add(2) <= WAD2_ipd;
	write_add(1) <= WAD1_ipd;
	write_add(0) <= WAD0_ipd;
      end if;

   end process;

   wrapper_write_data : process(WEN_ipd, WDATA3_ipd, WDATA2_ipd, WDATA1_ipd, WDATA0_ipd)

   begin
    if (WEN_ipd = '1') then
	DIN(3) <= WDATA3_ipd;
	DIN(2) <= WDATA2_ipd;
	DIN(1) <= WDATA1_ipd;
	DIN(0) <= WDATA0_ipd;
    else
	DIN <= x_data;
    end if;

   end process;


  VITALBehavior : PROCESS ( WEN_ipd, REN_ipd, WR_CLK, DIN, RD_ADD, WR_ADD)--, write_add)


   -- Temporary variables
   VARIABLE tempaddr 		: integer := 0;
   VARIABLE rd_address 		: integer := 0;
   VARIABLE rd_viol_flag 	: X01 := '0';

   -- Timing Check results
   VARIABLE Pviol_WCLK			: std_logic := '0';
   VARIABLE PeriodData_WCLK		: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_WR_ADD_stp_hld_0	: std_logic := '0';
   VARIABLE TimingData_WR_ADD_stp_hld_0	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_WR_ADD_stp_hld_1	: std_logic := '0';
   VARIABLE TimingData_WR_ADD_stp_hld_1	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_WR_ADD_stp_hld_2	: std_logic := '0';
   VARIABLE TimingData_WR_ADD_stp_hld_2	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_WR_ADD_stp_hld_3	: std_logic := '0';
   VARIABLE TimingData_WR_ADD_stp_hld_3	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_WR_ADD_stp_hld_4	: std_logic := '0';
   VARIABLE TimingData_WR_ADD_stp_hld_4	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_WR_DATA_stp_0		: std_logic := '0';
   VARIABLE TimingData_WR_DATA_stp_0	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_WR_DATA_stp_1		: std_logic := '0';
   VARIABLE TimingData_WR_DATA_stp_1	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_WR_DATA_stp_2		: std_logic := '0';
   VARIABLE TimingData_WR_DATA_stp_2	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_WR_DATA_stp_3		: std_logic := '0';
   VARIABLE TimingData_WR_DATA_stp_3	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_WEN_hld		: std_logic := '0';
   VARIABLE TimingData_WEN_hld		: VitalTimingDataType := VitalTimingDataInit;



 BEGIN
    -------------------------------------------------------------------
    -- Timing Check Section
    -------------------------------------------------------------------
    IF (TimingChecksOn) THEN


	VitalPeriodPulseCheck  (Pviol_WCLK,
				PeriodData_WCLK,
				WR_CLK, "WCLK",
				0.0 ns,
				0.0 ns,
				tpw_WCLK_posedge,
				0.0 ns,
				TRUE,
				InstancePath & "/RB_SA",
				TRUE,
				TRUE,
				WARNING );

	VitalSetupHoldCheck    (Tviol_WR_ADD_stp_hld_0,
				TimingData_WR_ADD_stp_hld_0,
				WR_ADD(0), "WAD0",
				0.0 ns,
				WR_CLK, "WCLK",
				0.0 ns,
				tsetup_WAD0_WCLK_noedge_posedge, tsetup_WAD0_WCLK_noedge_posedge, 
				thold_WAD0_WCLK_noedge_posedge, thold_WAD0_WCLK_noedge_posedge,
				TRUE,
				'/',
				InstancePath & "/RB_SA",
				TRUE,
				TRUE,
				WARNING );

	VitalSetupHoldCheck    (Tviol_WR_ADD_stp_hld_1,
				TimingData_WR_ADD_stp_hld_1,
				WR_ADD(1), "WAD1",
				0.0 ns,
				WR_CLK, "WCLK",
				0.0 ns,
				tsetup_WAD1_WCLK_noedge_posedge, tsetup_WAD1_WCLK_noedge_posedge, 
				thold_WAD1_WCLK_noedge_posedge, thold_WAD1_WCLK_noedge_posedge,
				TRUE,
				'/',
				InstancePath & "/RB_SA",
				TRUE,
				TRUE,
				WARNING );

	VitalSetupHoldCheck    (Tviol_WR_ADD_stp_hld_2,
				TimingData_WR_ADD_stp_hld_2,
				WR_ADD(2), "WAD2",
				0.0 ns,
				WR_CLK, "WCLK",
				0.0 ns,
				tsetup_WAD2_WCLK_noedge_posedge, tsetup_WAD2_WCLK_noedge_posedge, 
				thold_WAD2_WCLK_noedge_posedge, thold_WAD2_WCLK_noedge_posedge,
				TRUE,
				'/',
				InstancePath & "/RB_SA",
				TRUE,
				TRUE,
				WARNING );

	VitalSetupHoldCheck    (Tviol_WR_ADD_stp_hld_3,
				TimingData_WR_ADD_stp_hld_3,
				WR_ADD(3), "WAD3",
				0.0 ns,
				WR_CLK, "WCLK",
				0.0 ns,
				tsetup_WAD3_WCLK_noedge_posedge, tsetup_WAD3_WCLK_noedge_posedge, 
				thold_WAD3_WCLK_noedge_posedge, thold_WAD3_WCLK_noedge_posedge,
				TRUE,
				'/',
				InstancePath & "/RB_SA",
				TRUE,
				TRUE,
				WARNING );

	VitalSetupHoldCheck    (Tviol_WR_ADD_stp_hld_4,
				TimingData_WR_ADD_stp_hld_4,
				WR_ADD(4), "WAD4",
				0.0 ns,
				WR_CLK, "WCLK",
				0.0 ns,
				tsetup_WAD4_WCLK_noedge_posedge, tsetup_WAD4_WCLK_noedge_posedge, 
				thold_WAD4_WCLK_noedge_posedge, thold_WAD4_WCLK_noedge_posedge,
				TRUE,
				'/',
				InstancePath & "/RB_SA",
				TRUE,
				TRUE,
				WARNING );

	VitalSetupHoldCheck    (Tviol_WR_DATA_stp_0,
				TimingData_WR_DATA_stp_0,
				DIN(0), "WDATA0",
				0.0 ns,
				WR_CLK, "WCLK",
				0.0 ns,
				tsetup_WDATA0_WCLK_noedge_posedge, tsetup_WDATA0_WCLK_noedge_posedge, 
				thold_WDATA0_WCLK_noedge_posedge, thold_WDATA0_WCLK_noedge_posedge,
				TRUE,
				'/',
				InstancePath & "/RB_SA",
				TRUE,
				TRUE,
				WARNING );

	VitalSetupHoldCheck    (Tviol_WR_DATA_stp_1,
				TimingData_WR_DATA_stp_1,
				DIN(1), "WDATA1",
				0.0 ns,
				WR_CLK, "WCLK",
				0.0 ns,
				tsetup_WDATA1_WCLK_noedge_posedge, tsetup_WDATA1_WCLK_noedge_posedge, 
				thold_WDATA1_WCLK_noedge_posedge, thold_WDATA1_WCLK_noedge_posedge,
				TRUE,
				'/',
				InstancePath & "/RB_SA",
				TRUE,
				TRUE,
				WARNING );

	VitalSetupHoldCheck    (Tviol_WR_DATA_stp_2,
				TimingData_WR_DATA_stp_2,
				DIN(2), "WDATA2",
				0.0 ns,
				WR_CLK, "WCLK",
				0.0 ns,
				tsetup_WDATA2_WCLK_noedge_posedge, tsetup_WDATA2_WCLK_noedge_posedge, 
				thold_WDATA2_WCLK_noedge_posedge, thold_WDATA2_WCLK_noedge_posedge,
				TRUE,
				'/',
				InstancePath & "/RB_SA",
				TRUE,
				TRUE,
				WARNING );

	VitalSetupHoldCheck    (Tviol_WR_DATA_stp_3,
				TimingData_WR_DATA_stp_3,
				DIN(3), "WDATA3",
				0.0 ns,
				WR_CLK, "WCLK",
				0.0 ns,
				tsetup_WDATA3_WCLK_noedge_posedge, tsetup_WDATA3_WCLK_noedge_posedge, 
				thold_WDATA3_WCLK_noedge_posedge, thold_WDATA3_WCLK_noedge_posedge,
				TRUE,
				'/',
				InstancePath & "/RB_SA",
				TRUE,
				TRUE,
				WARNING );


	VitalSetupHoldCheck    (Tviol_WEN_hld,
				TimingData_WEN_hld,
				WEN_ipd, "WEN",
				0.0 ns,
				WR_CLK, "WCLK",
				0.0 ns,
				tsetup_WEN_WCLK_noedge_posedge,tsetup_WEN_WCLK_noedge_posedge,
				thold_WEN_WCLK_noedge_posedge,thold_WEN_WCLK_noedge_posedge,
				True,
				'/',
				InstancePath & "/RB_SA",
				TRUE,
				TRUE,
				WARNING );


    END IF; -- Timing Check Section


    -------------------------------------------------------------------
    -- Functionality Section
    -------------------------------------------------------------------

-- WRITE ADDRESS GOES XX

    if ( WR_CLK'EVENT and WR_CLK = '1' and vecX(WR_ADD)) then

        assert false
        report "Illegal Address Input: Undefined  Address at the Read_Write Port."
        severity note ;
        memory_array <= (others => x_data);

    end if;

-- ADDRESS HOLD AND SETUP VIOLATION EFFECT

    if( Tviol_WR_ADD_stp_hld_0 = 'X' or Tviol_WR_ADD_stp_hld_1 = 'X' or Tviol_WR_ADD_stp_hld_2 = 'X' or Tviol_WR_ADD_stp_hld_3 = 'X' or Tviol_WR_ADD_stp_hld_4 = 'X' ) then

        memory_array <= (others => x_data);

    else

-- DATA SETUP AND HOLD VIOLATION EFFECT

    if( Pviol_WCLK = 'X' or Tviol_WR_DATA_stp_0 = 'X' or Tviol_WR_DATA_stp_1 = 'X' or Tviol_WR_DATA_stp_2 = 'X' or Tviol_WR_DATA_stp_3 = 'X' or Tviol_WEN_hld = 'X') then
	tempaddr := vec2int(write_add);
	memory_array(tempaddr) <= x_data;
    end if;

    end if;

-- VALID MEMORY WRITE

    if ( WR_CLK'EVENT and WR_CLK = '1' and not(vecX(WR_ADD)) and not(Tviol_WR_ADD_stp_hld_0 = 'X' or Tviol_WR_ADD_stp_hld_1 = 'X' or Tviol_WR_ADD_stp_hld_2 = 'X' or Tviol_WR_ADD_stp_hld_3 = 'X' or Tviol_WR_ADD_stp_hld_4 = 'X') and not( Pviol_WCLK = 'X' or Tviol_WR_DATA_stp_0 = 'X' or Tviol_WR_DATA_stp_1 = 'X' or Tviol_WR_DATA_stp_2 = 'X' or Tviol_WR_DATA_stp_3 = 'X' or Tviol_WEN_hld = 'X') ) then
	tempaddr := vec2int(WR_ADD);
	memory_array(tempaddr) <= DIN;
    end if;

    if WR_CLK'EVENT and WR_CLK /= WCLK_ipd and WR_CLK'LAST_VALUE = '1' then
	memory_array(tempaddr) <= x_data;
    end if;


-- READ CYCLE VIOLATION EFFECT

    if(RD_ADD'EVENT  and REN_ipd = '1'  and vecX(RD_ADD)) then
	data_out <= x_data;
    elsif

-- VALID MEMORY READ


     (RD_ADD'EVENT  and REN_ipd = '1'  and not(vecX(RD_ADD))) then
	rd_address := vec2int(RD_ADD);
	data_out <= memory_array(rd_address);
    end if;


  END PROCESS;

    -------------------------------------------------------------------------------
    -- Temporary output signal should get assigned to the output signal.
    -------------------------------------------------------------------------------

  PROCESS(data_out, REN_ipd, RAD4_ipd, RAD3_ipd, RAD2_ipd, RAD1_ipd, RAD0_ipd) 

      VARIABLE RDATA3_1 : std_logic := 'X';
      VARIABLE RDATA2_1 : std_logic := 'X';
      VARIABLE RDATA1_1 : std_logic := 'X';
      VARIABLE RDATA0_1 : std_logic := 'X';
      VARIABLE GLITCH_DATA : VitalGlitchDataType;

   BEGIN
   
    RDATA0_1 := VitalBUF(data_out(0));    --- Is this Vital level0 compliant
    RDATA1_1 := VitalBUF(data_out(1));
    RDATA2_1 := VitalBUF(data_out(2));
    RDATA3_1 := VitalBUF(data_out(3));

      VitalPathDelay01 ( RDATA3, GLITCH_DATA, "RDATA3", RDATA3_1,
        Paths => (
        0 => ( REN_ipd'LAST_EVENT, tpd_REN_RDATA3, TRUE ),
        1 => ( RAD0_ipd'LAST_EVENT, tpd_RAD0_RDATA3, TRUE),
        2 => ( RAD1_ipd'LAST_EVENT, tpd_RAD1_RDATA3, TRUE),
        3 => ( RAD2_ipd'LAST_EVENT, tpd_RAD2_RDATA3, TRUE),
        4 => ( RAD3_ipd'LAST_EVENT, tpd_RAD3_RDATA3, TRUE),
        5 => ( RAD4_ipd'LAST_EVENT, tpd_RAD4_RDATA3, TRUE)),
        DefaultDelay=>VitalZeroDelay01,
        Mode=>VitalInertial,
        XON=>TRUE,
        MsgOn=>TRUE,
        MsgSeverity=>WARNING );

      VitalPathDelay01 ( RDATA2, GLITCH_DATA, "RDATA2", RDATA2_1,
        Paths => (
        0 => ( REN_ipd'LAST_EVENT, tpd_REN_RDATA2, TRUE ),
        1 => ( RAD0_ipd'LAST_EVENT, tpd_RAD0_RDATA2, TRUE),
        2 => ( RAD1_ipd'LAST_EVENT, tpd_RAD1_RDATA2, TRUE),
        3 => ( RAD2_ipd'LAST_EVENT, tpd_RAD2_RDATA2, TRUE),
        4 => ( RAD3_ipd'LAST_EVENT, tpd_RAD3_RDATA2, TRUE),
        5 => ( RAD4_ipd'LAST_EVENT, tpd_RAD4_RDATA2, TRUE)),
        DefaultDelay=>VitalZeroDelay01,
        Mode=>VitalInertial,
        XON=>TRUE,
        MsgOn=>TRUE,
        MsgSeverity=>WARNING );

      VitalPathDelay01 ( RDATA1, GLITCH_DATA, "RDATA1", RDATA1_1,
        Paths => (
        0 => ( REN_ipd'LAST_EVENT, tpd_REN_RDATA1, TRUE ),
        1 => ( RAD0_ipd'LAST_EVENT, tpd_RAD0_RDATA1, TRUE),
        2 => ( RAD1_ipd'LAST_EVENT, tpd_RAD1_RDATA1, TRUE),
        3 => ( RAD2_ipd'LAST_EVENT, tpd_RAD2_RDATA1, TRUE),
        4 => ( RAD3_ipd'LAST_EVENT, tpd_RAD3_RDATA1, TRUE),
        5 => ( RAD4_ipd'LAST_EVENT, tpd_RAD4_RDATA1, TRUE)),
        DefaultDelay=>VitalZeroDelay01,
        Mode=>VitalInertial,
        XON=>TRUE,
        MsgOn=>TRUE,
        MsgSeverity=>WARNING );

      VitalPathDelay01 ( RDATA0, GLITCH_DATA, "RDATA0", RDATA0_1,
        Paths => (
        0 => ( REN_ipd'LAST_EVENT, tpd_REN_RDATA0, TRUE ),
        1 => ( RAD0_ipd'LAST_EVENT, tpd_RAD0_RDATA0, TRUE),
        2 => ( RAD1_ipd'LAST_EVENT, tpd_RAD1_RDATA0, TRUE),
        3 => ( RAD2_ipd'LAST_EVENT, tpd_RAD2_RDATA0, TRUE),
        4 => ( RAD3_ipd'LAST_EVENT, tpd_RAD3_RDATA0, TRUE),
        5 => ( RAD4_ipd'LAST_EVENT, tpd_RAD4_RDATA0, TRUE)),
        DefaultDelay=>VitalZeroDelay01,
        Mode=>VitalInertial,
        XON=>TRUE,
        MsgOn=>TRUE,
        MsgSeverity=>WARNING );


END PROCESS;

END VITAL_VF;
configuration CFG_RB_SA_VITAL of RB_SA is
        for VITAL_VF
        end for;
end CFG_RB_SA_VITAL;
-----------------------------------------------------------------------


-----------------------------------------------------------------------
-- VITAL model for RB_SS 30.10 technology
-----------------------------------------------------------------------

LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.VITAL_timing.all;
USE IEEE.VITAL_primitives.all;
LIBRARY VF1;
USE VF1.ALL;
USE VF1.RAMPACK.ALL;

-----------------------------------------------------------------------
-- ENTITY declaration
-----------------------------------------------------------------------

ENTITY RB_SS IS
  GENERIC (
	tipd_WEN		: VitalDelayType01			:= (0.0 ns, 0.0 ns);
	tipd_REN		: VitalDelayType01			:= (0.0 ns, 0.0 ns);
	tipd_WCLK		: VitalDelayType01			:= (0.0 ns, 0.0 ns);
	tipd_RCLK		: VitalDelayType01			:= (0.0 ns, 0.0 ns);
	tipd_WDATA3		: VitalDelayType01 	   		:= (0.0 ns, 0.0 ns);
	tipd_WDATA2		: VitalDelayType01 	   		:= (0.0 ns, 0.0 ns);
	tipd_WDATA1		: VitalDelayType01 	   		:= (0.0 ns, 0.0 ns);
	tipd_WDATA0		: VitalDelayType01 	   		:= (0.0 ns, 0.0 ns);
	tipd_RAD4		: VitalDelayType01			:= (0.0 ns, 0.0 ns);
	tipd_RAD3		: VitalDelayType01			:= (0.0 ns, 0.0 ns);
	tipd_RAD2		: VitalDelayType01			:= (0.0 ns, 0.0 ns);
	tipd_RAD1		: VitalDelayType01			:= (0.0 ns, 0.0 ns);
	tipd_RAD0		: VitalDelayType01			:= (0.0 ns, 0.0 ns);
	tipd_WAD4		: VitalDelayType01			:= (0.0 ns, 0.0 ns);
	tipd_WAD3		: VitalDelayType01			:= (0.0 ns, 0.0 ns);
	tipd_WAD2		: VitalDelayType01			:= (0.0 ns, 0.0 ns);
	tipd_WAD1		: VitalDelayType01			:= (0.0 ns, 0.0 ns);
	tipd_WAD0		: VitalDelayType01			:= (0.0 ns, 0.0 ns);

	tsetup_WDATA3_WCLK_noedge_posedge		: VitalDelayType := 1.0 ns;
	tsetup_WDATA2_WCLK_noedge_posedge		: VitalDelayType := 1.0 ns;
	tsetup_WDATA1_WCLK_noedge_posedge		: VitalDelayType := 1.0 ns;
	tsetup_WDATA0_WCLK_noedge_posedge		: VitalDelayType := 1.0 ns;
	thold_WDATA3_WCLK_noedge_posedge		: VitalDelayType := 1.0 ns;
	thold_WDATA2_WCLK_noedge_posedge		: VitalDelayType := 1.0 ns;
	thold_WDATA1_WCLK_noedge_posedge		: VitalDelayType := 1.0 ns;
	thold_WDATA0_WCLK_noedge_posedge		: VitalDelayType := 1.0 ns;
	tsetup_WAD4_WCLK_noedge_posedge		: VitalDelayType := 1.0 ns;
	tsetup_WAD3_WCLK_noedge_posedge		: VitalDelayType := 1.0 ns;
	tsetup_WAD2_WCLK_noedge_posedge		: VitalDelayType := 1.0 ns;
	tsetup_WAD1_WCLK_noedge_posedge		: VitalDelayType := 1.0 ns;
	tsetup_WAD0_WCLK_noedge_posedge		: VitalDelayType := 1.0 ns;
	thold_WAD4_WCLK_noedge_posedge			: VitalDelayType := 1.0 ns;
	thold_WAD3_WCLK_noedge_posedge			: VitalDelayType := 1.0 ns;
	thold_WAD2_WCLK_noedge_posedge			: VitalDelayType := 1.0 ns;
	thold_WAD1_WCLK_noedge_posedge			: VitalDelayType := 1.0 ns;
	thold_WAD0_WCLK_noedge_posedge			: VitalDelayType := 1.0 ns;
	tpw_WCLK_posedge					: VitalDelayType := 1.0 ns;
	tsetup_WEN_WCLK_noedge_posedge			: VitalDelayType := 1.0 ns;
	thold_WEN_WCLK_noedge_posedge			: VitalDelayType := 1.0 ns;
	tsetup_RAD4_RCLK_noedge_posedge		: VitalDelayType := 1.0 ns;
	tsetup_RAD3_RCLK_noedge_posedge		: VitalDelayType := 1.0 ns;
	tsetup_RAD2_RCLK_noedge_posedge		: VitalDelayType := 1.0 ns;
	tsetup_RAD1_RCLK_noedge_posedge		: VitalDelayType := 1.0 ns;
	tsetup_RAD0_RCLK_noedge_posedge		: VitalDelayType := 1.0 ns;
	thold_RAD4_RCLK_noedge_posedge			: VitalDelayType := 1.0 ns;
	thold_RAD3_RCLK_noedge_posedge			: VitalDelayType := 1.0 ns;
	thold_RAD2_RCLK_noedge_posedge			: VitalDelayType := 1.0 ns;
	thold_RAD1_RCLK_noedge_posedge			: VitalDelayType := 1.0 ns;
	thold_RAD0_RCLK_noedge_posedge			: VitalDelayType := 1.0 ns;
	tpd_RCLK_RDATA3				: VitalDelayType01 := (2.0 ns,2.0 ns);
	tpd_RCLK_RDATA2				: VitalDelayType01 := (2.0 ns,2.0 ns);
	tpd_RCLK_RDATA1				: VitalDelayType01 := (2.0 ns,2.0 ns);
	tpd_RCLK_RDATA0				: VitalDelayType01 := (2.0 ns,2.0 ns);
	tpw_RCLK_posedge				: VitalDelayType := 1.0 ns;
	tsetup_REN_RCLK_noedge_posedge			: VitalDelayType := 1.0 ns;
	thold_REN_RCLK_noedge_posedge			: VitalDelayType := 1.0 ns;

	TimingChecksOn : BOOLEAN := TRUE;
	MsgOn : BOOLEAN := TRUE;
	XON : BOOLEAN := TRUE;
	InstancePath : STRING := "*"
            );
  PORT	(
	WEN		: IN	std_logic ;
	REN		: IN	std_logic ;
	RDATA3		: OUT	std_logic ;
	RDATA2		: OUT	std_logic ;
	RDATA1		: OUT	std_logic ;
	RDATA0		: OUT	std_logic ;
	WCLK		: IN	std_logic ;
	RCLK		: IN	std_logic ;
	WDATA3	        : IN	std_logic ;
	WDATA2	        : IN	std_logic ;
	WDATA1	        : IN	std_logic ;
	WDATA0	        : IN	std_logic ;
	RAD4		: IN	std_logic ;
	RAD3		: IN	std_logic ;
	RAD2		: IN	std_logic ;
	RAD1		: IN	std_logic ;
	RAD0		: IN	std_logic ;
	WAD4		: IN	std_logic ;
	WAD3		: IN	std_logic ;
	WAD2		: IN	std_logic ;
	WAD1		: IN	std_logic ;
	WAD0		: IN	std_logic
	);


   ATTRIBUTE VITAL_LEVEL0 OF RB_SS : ENTITY IS TRUE;

END RB_SS;

-----------------------------------------------------------------------
-- ARCHITECTURE declaration
-----------------------------------------------------------------------
ARCHITECTURE VITAL_VF OF RB_SS IS

    ATTRIBUTE VITAL_LEVEL1 OF VITAL_VF : ARCHITECTURE IS FALSE;

	SIGNAL WEN_ipd		: std_logic := 'X'; 
	SIGNAL REN_ipd		: std_logic := 'X';
	SIGNAL WCLK_ipd		: std_logic := '0';
	SIGNAL WR_CLK		: std_logic := '0';
	SIGNAL RCLK_ipd		: std_logic := '0';
	SIGNAL RD_CLK		: std_logic := '0';
	SIGNAL WDATA3_ipd	: std_logic := '0';
	SIGNAL WDATA2_ipd	: std_logic := '0';
	SIGNAL WDATA1_ipd	: std_logic := '0';
	SIGNAL WDATA0_ipd	: std_logic := '0';
	SIGNAL DIN		: std_logic_vector(3 DOWNTO 0);
	SIGNAL RAD4_ipd		: std_logic := '0';
	SIGNAL RAD3_ipd		: std_logic := '0';
	SIGNAL RAD2_ipd		: std_logic := '0';
	SIGNAL RAD1_ipd		: std_logic := '0';
	SIGNAL RAD0_ipd		: std_logic := '0';
	SIGNAL RD_ADD		: std_logic_vector(4 DOWNTO 0);
	SIGNAL WAD4_ipd		: std_logic := '0';
	SIGNAL WAD3_ipd		: std_logic := '0';
	SIGNAL WAD2_ipd		: std_logic := '0';
	SIGNAL WAD1_ipd		: std_logic := '0';
	SIGNAL WAD0_ipd		: std_logic := '0';
	SIGNAL WR_ADD		: std_logic_vector(4 DOWNTO 0);
	SIGNAL write_add	: std_logic_vector(4 DOWNTO 0);
	SIGNAL data_out		: std_logic_vector(3 DOWNTO 0);
	--SIGNAL output_delay	: time		:= 0 ns;

BEGIN
   
  ---------------------------------------------------------------------
  -- INPUT PATH DELAYs
  ---------------------------------------------------------------------
  WIREDELAY : BLOCK
  BEGIN
	VitalWireDelay (WEN_ipd,		WEN,		tipd_WEN);
	VitalWireDelay (REN_ipd,		REN,		tipd_REN);
	VitalWireDelay (WCLK_ipd,		WCLK,		tipd_WCLK);
	VitalWireDelay (RCLK_ipd,		RCLK,		tipd_RCLK);
	VitalWireDelay (WDATA0_ipd,		WDATA0,		tipd_WDATA0);
	VitalWireDelay (WDATA1_ipd,		WDATA1,		tipd_WDATA1);
	VitalWireDelay (WDATA2_ipd,		WDATA2,		tipd_WDATA2);
	VitalWireDelay (WDATA3_ipd,		WDATA3,		tipd_WDATA3);
	VitalWireDelay (RAD0_ipd,		RAD0,		tipd_RAD0);
	VitalWireDelay (RAD1_ipd,		RAD1,		tipd_RAD1);
	VitalWireDelay (RAD2_ipd,		RAD2,		tipd_RAD2);
	VitalWireDelay (RAD3_ipd,		RAD3,		tipd_RAD3);
	VitalWireDelay (RAD4_ipd,		RAD4,		tipd_RAD4);
	VitalWireDelay (WAD0_ipd,		WAD0,		tipd_WAD0);
	VitalWireDelay (WAD1_ipd,		WAD1,		tipd_WAD1);
	VitalWireDelay (WAD2_ipd,		WAD2,		tipd_WAD2);
	VitalWireDelay (WAD3_ipd,		WAD3,		tipd_WAD3);
	VitalWireDelay (WAD4_ipd,		WAD4,		tipd_WAD4);

  END BLOCK;

  ---------------------------------------------------------------------
  -- Behavior Section
  ---------------------------------------------------------------------

  ---------------------------------------------------------------------
  -- Wrapper Section
  ---------------------------------------------------------------------

   wrapper_read_add : process(REN_ipd, RAD4_ipd, RAD3_ipd, RAD2_ipd, RAD1_ipd, RAD0_ipd)

   begin
    if (REN_ipd = '1') then
	RD_ADD(0) <= RAD0_ipd;
	RD_ADD(1) <= RAD1_ipd;
	RD_ADD(2) <= RAD2_ipd;
	RD_ADD(3) <= RAD3_ipd;
	RD_ADD(4) <= RAD4_ipd;
    else
	RD_ADD <= x_add;
    end if;

   end process;

   wrapper_read_clk : process(REN_ipd, RCLK_ipd)

   begin
    if (REN_ipd = '1') then
	RD_CLK <= RCLK_ipd;
    else
	RD_CLK <= '0';
    end if;

   end process;

   wrapper_write_add : process(WEN_ipd, WAD4_ipd, WAD3_ipd, WAD2_ipd, WAD1_ipd, WAD0_ipd)

   begin
--   if (WEN_ipd = '1') then
	WR_ADD(0) <= WAD0_ipd;
	WR_ADD(1) <= WAD1_ipd;
	WR_ADD(2) <= WAD2_ipd;
	WR_ADD(3) <= WAD3_ipd;
	WR_ADD(4) <= WAD4_ipd;
 --   else
--	WR_ADD <= x_add;
 --  end if;

   end process;

   wrapper_write_clk : process(WEN_ipd, WCLK_ipd)

   begin
    if (WEN_ipd = '1') then
	WR_CLK <= WCLK_ipd;
    else
	WR_CLK <= '0';
    end if;

   end process;

   process(WR_CLK)

    begin
      if WR_CLK = '1' then
	write_add(0) <= WAD0_ipd;
	write_add(1) <= WAD1_ipd;
	write_add(2) <= WAD2_ipd;
	write_add(3) <= WAD3_ipd;
	write_add(4) <= WAD4_ipd;
      end if;

   end process;

   wrapper_write_data : process(WEN_ipd, WDATA3_ipd,WDATA2_ipd, WDATA1_ipd, WDATA0_ipd)

   begin
    if (WEN_ipd = '1') then
	DIN(0) <= WDATA0_ipd;
	DIN(1) <= WDATA1_ipd;
	DIN(2) <= WDATA2_ipd;
	DIN(3) <= WDATA3_ipd;
    else
	DIN <= x_data;
    end if;

   end process;


  VITALBehavior : PROCESS ( WEN_ipd, REN_ipd, WR_CLK, RD_CLK, DIN, RD_ADD, WR_ADD )

   VARIABLE memory_array : memory_array_typ;

   -- Temporary variables
   VARIABLE tempaddr : integer := 0;
   VARIABLE rd_address : integer := 0;

   -- Timing Check results
   VARIABLE Pviol_RCLK			: std_logic := '0';
   VARIABLE PeriodData_RCLK		: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_WCLK			: std_logic := '0';
   VARIABLE PeriodData_WCLK		: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_WR_ADD_stp_hld_0	: std_logic := '0';
   VARIABLE TimingData_WR_ADD_stp_hld_0	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_WR_ADD_stp_hld_1	: std_logic := '0';
   VARIABLE TimingData_WR_ADD_stp_hld_1	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_WR_ADD_stp_hld_2	: std_logic := '0';
   VARIABLE TimingData_WR_ADD_stp_hld_2	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_WR_ADD_stp_hld_3	: std_logic := '0';
   VARIABLE TimingData_WR_ADD_stp_hld_3	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_WR_ADD_stp_hld_4	: std_logic := '0';
   VARIABLE TimingData_WR_ADD_stp_hld_4	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_WR_DATA_stp_0		: std_logic := '0';
   VARIABLE TimingData_WR_DATA_stp_0	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_WR_DATA_stp_1		: std_logic := '0';
   VARIABLE TimingData_WR_DATA_stp_1	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_WR_DATA_stp_2		: std_logic := '0';
   VARIABLE TimingData_WR_DATA_stp_2	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_WR_DATA_stp_3		: std_logic := '0';
   VARIABLE TimingData_WR_DATA_stp_3	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_WR_DATA_hld_0		: std_logic := '0';
   VARIABLE TimingData_WR_DATA_hld_0	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_WR_DATA_hld_1		: std_logic := '0';
   VARIABLE TimingData_WR_DATA_hld_1	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_WR_DATA_hld_2		: std_logic := '0';
   VARIABLE TimingData_WR_DATA_hld_2	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_WR_DATA_hld_3		: std_logic := '0';
   VARIABLE TimingData_WR_DATA_hld_3	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_RD_ADD_stp_hld_0	: std_logic := '0';
   VARIABLE TimingData_RD_ADD_stp_hld_0	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_RD_ADD_stp_hld_1	: std_logic := '0';
   VARIABLE TimingData_RD_ADD_stp_hld_1	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_RD_ADD_stp_hld_2	: std_logic := '0';
   VARIABLE TimingData_RD_ADD_stp_hld_2	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_RD_ADD_stp_hld_3	: std_logic := '0';
   VARIABLE TimingData_RD_ADD_stp_hld_3	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_RD_ADD_stp_hld_4	: std_logic := '0';
   VARIABLE TimingData_RD_ADD_stp_hld_4	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_WEN_hld		: std_logic := '0';
   VARIABLE TimingData_WEN_hld		: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_REN_hld		: std_logic := '0';
   VARIABLE TimingData_REN_hld		: VitalTimingDataType := VitalTimingDataInit;



 BEGIN
    -------------------------------------------------------------------
    -- Timing Check Section
    -------------------------------------------------------------------
    IF (TimingChecksOn) THEN

	VitalPeriodPulseCheck  (Pviol_RCLK,
				PeriodData_RCLK,
				RD_CLK, "RCLK",
				0.0 ns,
				0.0 ns,
				tpw_RCLK_posedge,
				0.0 ns,
				TRUE,
				InstancePath & "/RB_SS",
				TRUE,
				TRUE,
				WARNING );

	VitalPeriodPulseCheck  (Pviol_WCLK,
				PeriodData_WCLK,
				WR_CLK, "WCLK",
				0.0 ns,
				0.0 ns,
				tpw_WCLK_posedge,
				0.0 ns,
				TRUE,
				InstancePath & "/RB_SS",
				TRUE,
				TRUE,
				WARNING );

	VitalSetupHoldCheck    (Tviol_WR_ADD_stp_hld_0,
				TimingData_WR_ADD_stp_hld_0,
				WR_ADD(0), "WAD0",
				0.0 ns,
				WR_CLK, "WCLK",
				0.0 ns,
				tsetup_WAD0_WCLK_noedge_posedge, tsetup_WAD0_WCLK_noedge_posedge, 
				thold_WAD0_WCLK_noedge_posedge, thold_WAD0_WCLK_noedge_posedge,
				WEN_ipd = '1',
				'/',
				InstancePath & "/RB_SS",
				TRUE,
				TRUE,
				WARNING );

	VitalSetupHoldCheck    (Tviol_WR_ADD_stp_hld_1,
				TimingData_WR_ADD_stp_hld_1,
				WR_ADD(1), "WAD1",
				0.0 ns,
				WR_CLK, "WCLK",
				0.0 ns,
				tsetup_WAD1_WCLK_noedge_posedge, tsetup_WAD1_WCLK_noedge_posedge, 
				thold_WAD1_WCLK_noedge_posedge, thold_WAD1_WCLK_noedge_posedge,
				WEN_ipd = '1',
				'/',
				InstancePath & "/RB_SS",
				TRUE,
				TRUE,
				WARNING );

	VitalSetupHoldCheck    (Tviol_WR_ADD_stp_hld_2,
				TimingData_WR_ADD_stp_hld_2,
				WR_ADD(2), "WAD2",
				0.0 ns,
				WR_CLK, "WCLK",
				0.0 ns,
				tsetup_WAD2_WCLK_noedge_posedge, tsetup_WAD2_WCLK_noedge_posedge, 
				thold_WAD2_WCLK_noedge_posedge, thold_WAD2_WCLK_noedge_posedge,
				WEN_ipd = '1',
				'/',
				InstancePath & "/RB_SS",
				TRUE,
				TRUE,
				WARNING );

	VitalSetupHoldCheck    (Tviol_WR_ADD_stp_hld_3,
				TimingData_WR_ADD_stp_hld_3,
				WR_ADD(3), "WAD3",
				0.0 ns,
				WR_CLK, "WCLK",
				0.0 ns,
				tsetup_WAD3_WCLK_noedge_posedge, tsetup_WAD3_WCLK_noedge_posedge, 
				thold_WAD3_WCLK_noedge_posedge, thold_WAD3_WCLK_noedge_posedge,
				WEN_ipd = '1',
				'/',
				InstancePath & "/RB_SS",
				TRUE,
				TRUE,
				WARNING );

	VitalSetupHoldCheck    (Tviol_WR_ADD_stp_hld_4,
				TimingData_WR_ADD_stp_hld_4,
				WR_ADD(4), "WAD4",
				0.0 ns,
				WR_CLK, "WCLK",
				0.0 ns,
				tsetup_WAD4_WCLK_noedge_posedge, tsetup_WAD4_WCLK_noedge_posedge, 
				thold_WAD4_WCLK_noedge_posedge, thold_WAD4_WCLK_noedge_posedge,
				WEN_ipd = '1',
				'/',
				InstancePath & "/RB_SS",
				TRUE,
				TRUE,
				WARNING );

	VitalSetupHoldCheck    (Tviol_WR_DATA_stp_0,
				TimingData_WR_DATA_stp_0,
				DIN(0), "WDATA0",
				0.0 ns,
				WR_CLK, "WCLK",
				0.0 ns,
				tsetup_WDATA0_WCLK_noedge_posedge, tsetup_WDATA0_WCLK_noedge_posedge, 
				0.0 ns, 0.0 ns,
				WEN_ipd = '1',
				'/',
				InstancePath & "/RB_SS",
				TRUE,
				TRUE,
				WARNING );

	VitalSetupHoldCheck    (Tviol_WR_DATA_stp_1,
				TimingData_WR_DATA_stp_1,
				DIN(1), "WDATA1",
				0.0 ns,
				WR_CLK, "WCLK",
				0.0 ns,
				tsetup_WDATA1_WCLK_noedge_posedge, tsetup_WDATA1_WCLK_noedge_posedge, 
				0.0 ns, 0.0 ns,
				WEN_ipd = '1',
				'/',
				InstancePath & "/RB_SS",
				TRUE,
				TRUE,
				WARNING );

	VitalSetupHoldCheck    (Tviol_WR_DATA_stp_2,
				TimingData_WR_DATA_stp_2,
				DIN(2), "WDATA2",
				0.0 ns,
				WR_CLK, "WCLK",
				0.0 ns,
				tsetup_WDATA2_WCLK_noedge_posedge, tsetup_WDATA2_WCLK_noedge_posedge, 
				0.0 ns, 0.0 ns,
				WEN_ipd = '1',
				'/',
				InstancePath & "/RB_SS",
				TRUE,
				TRUE,
				WARNING );

	VitalSetupHoldCheck    (Tviol_WR_DATA_stp_3,
				TimingData_WR_DATA_stp_3,
				DIN(3), "WDATA3",
				0.0 ns,
				WR_CLK, "WCLK",
				0.0 ns,
				tsetup_WDATA3_WCLK_noedge_posedge, tsetup_WDATA3_WCLK_noedge_posedge, 
				0.0 ns, 0.0 ns,
				WEN_ipd = '1',
				'/',
				InstancePath & "/RB_SS",
				TRUE,
				TRUE,
				WARNING );

	VitalSetupHoldCheck    (Tviol_WR_DATA_hld_0,
				TimingData_WR_DATA_hld_0,
				DIN(0), "WDATA0",
				0.0 ns,
				WR_CLK, "WCLK",
				0.0 ns,
				0.0 ns, 0.0 ns,
				thold_WDATA0_WCLK_noedge_posedge, thold_WDATA0_WCLK_noedge_posedge,
				WEN_ipd = '1',
				'/',
				InstancePath & "/RB_SS",
				TRUE,
				TRUE,
				WARNING );

	VitalSetupHoldCheck    (Tviol_WR_DATA_hld_1,
				TimingData_WR_DATA_hld_1,
				DIN(1), "WDATA1",
				0.0 ns,
				WR_CLK, "WCLK",
				0.0 ns,
				0.0 ns, 0.0 ns,
				thold_WDATA1_WCLK_noedge_posedge, thold_WDATA1_WCLK_noedge_posedge,
				WEN_ipd = '1',
				'/',
				InstancePath & "/RB_SS",
				TRUE,
				TRUE,
				WARNING );

	VitalSetupHoldCheck    (Tviol_WR_DATA_hld_2,
				TimingData_WR_DATA_hld_2,
				DIN(2), "WDATA2",
				0.0 ns,
				WR_CLK, "WCLK",
				0.0 ns,
				0.0 ns, 0.0 ns,
				thold_WDATA2_WCLK_noedge_posedge, thold_WDATA2_WCLK_noedge_posedge,
				WEN_ipd = '1',
				'/',
				InstancePath & "/RB_SS",
				TRUE,
				TRUE,
				WARNING );

	VitalSetupHoldCheck    (Tviol_WR_DATA_hld_3,
				TimingData_WR_DATA_hld_3,
				DIN(3), "WDATA3",
				0.0 ns,
				WR_CLK, "WCLK",
				0.0 ns,
				0.0 ns, 0.0 ns,
				thold_WDATA3_WCLK_noedge_posedge, thold_WDATA3_WCLK_noedge_posedge,
				WEN_ipd = '1',
				'/',
				InstancePath & "/RB_SS",
				TRUE,
				TRUE,
				WARNING );

	VitalSetupHoldCheck    (Tviol_RD_ADD_stp_hld_0,
				TimingData_RD_ADD_stp_hld_0,
				RD_ADD(0), "RAD0",
				0.0 ns,
				RD_CLK, "RCLK",
				0.0 ns,
				tsetup_RAD0_RCLK_noedge_posedge, tsetup_RAD0_RCLK_noedge_posedge, 
				thold_RAD0_RCLK_noedge_posedge, thold_RAD0_RCLK_noedge_posedge,
				REN_ipd = '1',
				'/',
				InstancePath & "/RB_SS",
				TRUE,
				TRUE,
				WARNING );

	VitalSetupHoldCheck    (Tviol_RD_ADD_stp_hld_1,
				TimingData_RD_ADD_stp_hld_1,
				RD_ADD(1), "RAD1",
				0.0 ns,
				RD_CLK, "RCLK",
				0.0 ns,
				tsetup_RAD1_RCLK_noedge_posedge, tsetup_RAD1_RCLK_noedge_posedge, 
				thold_RAD1_RCLK_noedge_posedge, thold_RAD1_RCLK_noedge_posedge,
				REN_ipd = '1',
				'/',
				InstancePath & "/RB_SS",
				TRUE,
				TRUE,
				WARNING );

	VitalSetupHoldCheck    (Tviol_RD_ADD_stp_hld_2,
				TimingData_RD_ADD_stp_hld_2,
				RD_ADD(2), "RAD2",
				0.0 ns,
				RD_CLK, "RCLK",
				0.0 ns,
				tsetup_RAD2_RCLK_noedge_posedge, tsetup_RAD2_RCLK_noedge_posedge, 
				thold_RAD2_RCLK_noedge_posedge, thold_RAD2_RCLK_noedge_posedge,
				REN_ipd = '1',
				'/',
				InstancePath & "/RB_SS",
				TRUE,
				TRUE,
				WARNING );

	VitalSetupHoldCheck    (Tviol_RD_ADD_stp_hld_3,
				TimingData_RD_ADD_stp_hld_3,
				RD_ADD(3), "RAD3",
				0.0 ns,
				RD_CLK, "RCLK",
				0.0 ns,
				tsetup_RAD3_RCLK_noedge_posedge, tsetup_RAD3_RCLK_noedge_posedge, 
				thold_RAD3_RCLK_noedge_posedge, thold_RAD3_RCLK_noedge_posedge,
				REN_ipd = '1',
				'/',
				InstancePath & "/RB_SS",
				TRUE,
				TRUE,
				WARNING );

	VitalSetupHoldCheck    (Tviol_RD_ADD_stp_hld_4,
				TimingData_RD_ADD_stp_hld_4,
				RD_ADD(4), "RAD4",
				0.0 ns,
				RD_CLK, "RCLK",
				0.0 ns,
				tsetup_RAD4_RCLK_noedge_posedge, tsetup_RAD4_RCLK_noedge_posedge, 
				thold_RAD4_RCLK_noedge_posedge, thold_RAD4_RCLK_noedge_posedge,
				REN_ipd = '1',
				'/',
				InstancePath & "/RB_SS",
				TRUE,
				TRUE,
				WARNING );

	VitalSetupHoldCheck    (Tviol_WEN_hld,
				TimingData_WEN_hld,
				WEN_ipd, "WEN",
				0.0 ns,
				WR_CLK, "WCLK",
				0.0 ns,
				tsetup_WEN_WCLK_noedge_posedge,thold_WEN_WCLK_noedge_posedge,
				tsetup_WEN_WCLK_noedge_posedge,thold_WEN_WCLK_noedge_posedge,
				True,
				'/',
				InstancePath & "/RB_SS",
				TRUE,
				TRUE,
				WARNING );

	VitalSetupHoldCheck    (Tviol_REN_hld,
				TimingData_REN_hld,
				REN_ipd, "REN",
				0.0 ns,
				RD_CLK, "RCLK",
                                0.0 ns,
				tsetup_REN_RCLK_noedge_posedge,thold_REN_RCLK_noedge_posedge,
				tsetup_REN_RCLK_noedge_posedge,thold_REN_RCLK_noedge_posedge,
				True,
				'/',
				InstancePath & "/RB_SS",
				TRUE,
				TRUE,
				WARNING );

    END IF; -- Timing Check Section

    -------------------------------------------------------------------
    -- Functionality Section
    -------------------------------------------------------------------

-- WRITE ADDRESS GOES XX

    if ( WR_CLK'EVENT and WR_CLK = '1' and vecX(WR_ADD)) then

        assert false
        report "Illegal Address Input: Undefined  Address at the Write Port."
        severity note ;
        memory_array := (others => x_data);

    end if;

-- ADDRESS HOLD AND SETUP VIOLATION EFFECT

    if( Tviol_WR_ADD_stp_hld_0 = 'X' or Tviol_WR_ADD_stp_hld_1 = 'X' or Tviol_WR_ADD_stp_hld_2 = 'X' or Tviol_WR_ADD_stp_hld_3 = 'X' or Tviol_WR_ADD_stp_hld_4 = 'X' ) then

        memory_array := (others => x_data);

    else

-- DATA SETUP AND HOLD VIOLATION EFFECT

    if( Pviol_WCLK = 'X' or Tviol_WR_DATA_hld_0 = 'X' or Tviol_WR_DATA_hld_1 = 'X' or Tviol_WR_DATA_hld_2 = 'X' or Tviol_WR_DATA_hld_3 = 'X' or Tviol_WEN_hld = 'X') then
	tempaddr := vec2int(write_add);
	memory_array(tempaddr) := x_data;
    end if;

    if( Tviol_WR_DATA_stp_0 = 'X' or Tviol_WR_DATA_stp_1 = 'X' or Tviol_WR_DATA_stp_2 = 'X' or Tviol_WR_DATA_stp_3 = 'X') then
	tempaddr := vec2int(WR_ADD);
	memory_array(tempaddr) := x_data;
    end if;

    end if;

-- VALID MEMORY WRITE

    if ( WR_CLK'EVENT and WR_CLK = '1' and not(vecX(WR_ADD)) and not(Tviol_WR_ADD_stp_hld_0 = 'X' or Tviol_WR_ADD_stp_hld_1 = 'X' or Tviol_WR_ADD_stp_hld_2 = 'X' or Tviol_WR_ADD_stp_hld_3 = 'X' or Tviol_WR_ADD_stp_hld_4 = 'X') and not( Pviol_WCLK = 'X' or Tviol_WR_DATA_hld_0 = 'X' or Tviol_WR_DATA_hld_1 = 'X' or Tviol_WR_DATA_hld_2 = 'X' or Tviol_WR_DATA_hld_3 = 'X' or Tviol_WEN_hld = 'X') and not( Tviol_WR_DATA_stp_0 = 'X' or Tviol_WR_DATA_stp_1 = 'X' or Tviol_WR_DATA_stp_2 = 'X' or Tviol_WR_DATA_stp_3 = 'X')) then
	tempaddr := vec2int(WR_ADD);
	memory_array(tempaddr) := DIN;
    end if;

    if WR_CLK'EVENT and WR_CLK /= WCLK_ipd and WR_CLK'LAST_VALUE = '1' then
	memory_array(tempaddr) := x_data;
    end if;


-- READ ADDRESS CYCLE VIOLATION EFFECT

    if( Tviol_RD_ADD_stp_hld_0 = 'X' or Tviol_RD_ADD_stp_hld_1 = 'X' or Tviol_RD_ADD_stp_hld_2 = 'X' or Tviol_RD_ADD_stp_hld_3 = 'X' or Tviol_RD_ADD_stp_hld_4 = 'X' or Pviol_RCLK = 'X' or Tviol_REN_hld = 'X' or (RD_CLK'EVENT and RD_CLK = '1' and vecX(RD_ADD))) then
	--output_delay <= 0 ns;
	data_out <= x_data;
    elsif

-- VALID MEMORY READ

    (RD_CLK'EVENT and RD_CLK = '1' and not( Tviol_RD_ADD_stp_hld_0 = 'X' or Tviol_RD_ADD_stp_hld_1 = 'X' or Tviol_RD_ADD_stp_hld_2 = 'X' or Tviol_RD_ADD_stp_hld_3 = 'X' or Tviol_RD_ADD_stp_hld_4 = 'X' or Pviol_RCLK = 'X' or Tviol_REN_hld = 'X' or vecX(RD_ADD)) ) then
	rd_address := vec2int(RD_ADD);
	--output_delay <= tpd_RCLK_RDATA3_posedge;
	data_out <= memory_array(rd_address);
    end if;

    if RD_CLK'EVENT and RD_CLK /= RCLK_ipd and RD_CLK'LAST_VALUE = '1' then
	--output_delay <= 0 ns;
	data_out <= x_data;
    end if;


  END PROCESS;

    -------------------------------------------------------------------------------
    -- Temporary output signal should get assigned to the output signal.
    -------------------------------------------------------------------------------

  PROCESS(data_out, RCLK_ipd)

   VARIABLE RDATA0_1 : std_logic := 'X';
   VARIABLE RDATA1_1 : std_logic := 'X';
   VARIABLE RDATA2_1 : std_logic := 'X';
   VARIABLE RDATA3_1 : std_logic := 'X';
   VARIABLE GLITCH_DATA : VitalGlitchDataType;
  BEGIN

    RDATA0_1 := VitalBUF(data_out(0));    --- Is this Vital level0 compliant
    RDATA1_1 := VitalBUF(data_out(1)); 
    RDATA2_1 := VitalBUF(data_out(2)); 
    RDATA3_1 := VitalBUF(data_out(3)); 
    
      VitalPathDelay01 ( RDATA3, GLITCH_DATA, "RDATA3", RDATA3_1,
        Paths => (
        0 => ( RCLK_ipd'LAST_EVENT, tpd_RCLK_RDATA3, TRUE ) ),
        DefaultDelay=>VitalZeroDelay01,
        Mode=>VitalInertial,
        XON=>TRUE,
        MsgOn=>TRUE,
        MsgSeverity=>WARNING );
    
      VitalPathDelay01 ( RDATA2, GLITCH_DATA, "RDATA2", RDATA2_1,
        Paths => (
        0 => ( RCLK_ipd'LAST_EVENT, tpd_RCLK_RDATA2, TRUE ) ),
        DefaultDelay=>VitalZeroDelay01,
        Mode=>VitalInertial,
        XON=>TRUE,
        MsgOn=>TRUE,
        MsgSeverity=>WARNING );

      VitalPathDelay01 ( RDATA1, GLITCH_DATA, "RDATA1", RDATA1_1,
        Paths => (
        0 => ( RCLK_ipd'LAST_EVENT, tpd_RCLK_RDATA1, TRUE ) ),
        DefaultDelay=>VitalZeroDelay01,
        Mode=>VitalInertial,
        XON=>TRUE,
        MsgOn=>TRUE,
        MsgSeverity=>WARNING );

      VitalPathDelay01 ( RDATA0, GLITCH_DATA, "RDATA0", RDATA0_1,
        Paths => (
        0 => ( RCLK_ipd'LAST_EVENT, tpd_RCLK_RDATA0, TRUE ) ),
        DefaultDelay=>VitalZeroDelay01,
        Mode=>VitalInertial,
        XON=>TRUE,
        MsgOn=>TRUE,
        MsgSeverity=>WARNING );

END PROCESS;

END VITAL_VF;
configuration CFG_RB_SS_VITAL of RB_SS is
        for VITAL_VF
        end for;
end CFG_RB_SS_VITAL;
-------------------------------------------------------------------
-- VITAL model for RB_DAR 30.10 technology 
----------------------------------------------------------------------- 
 
LIBRARY IEEE; 
USE IEEE.std_logic_1164.ALL; 
USE IEEE.VITAL_timing.all; 
USE IEEE.std_logic_textio.all; 
USE IEEE.VITAL_primitives.all; 
LIBRARY std; 
USE std.textio.all; 
LIBRARY VF1; 
USE VF1.ALL; 
USE VF1.RAMPACK.ALL; 
 
----------------------------------------------------------------------- 
-- ENTITY declaration 
----------------------------------------------------------------------- 
 
ENTITY RB_DAR IS 
  GENERIC ( 
	tipd_WEN		: VitalDelayType01			:= (0.0 ns, 0.0 ns); 
	tipd_REN		: VitalDelayType01			:= (0.0 ns, 0.0 ns); 
	tipd_WRCLK		: VitalDelayType01			:= (0.0 ns, 0.0 ns); 
	tipd_ADRCLK		: VitalDelayType01			:= (0.0 ns, 0.0 ns); 
	tipd_OE		: VitalDelayType01			:= (0.0 ns, 0.0 ns); 
        tipd_WRDATA3            : VitalDelayType01      := (0.0 ns, 0.0 ns);
        tipd_WRDATA2            : VitalDelayType01      := (0.0 ns, 0.0 ns);
        tipd_WRDATA1            : VitalDelayType01      := (0.0 ns, 0.0 ns);
        tipd_WRDATA0            : VitalDelayType01      := (0.0 ns, 0.0 ns);
        tipd_WRAD4              : VitalDelayType01      := (0.0 ns, 0.0 ns);
        tipd_WRAD3              : VitalDelayType01      := (0.0 ns, 0.0 ns);
        tipd_WRAD2              : VitalDelayType01      := (0.0 ns, 0.0 ns);
        tipd_WRAD1              : VitalDelayType01      := (0.0 ns, 0.0 ns);
        tipd_WRAD0              : VitalDelayType01      := (0.0 ns, 0.0 ns);
        tipd_RAD4              : VitalDelayType01      := (0.0 ns, 0.0 ns);
        tipd_RAD3              : VitalDelayType01      := (0.0 ns, 0.0 ns);
        tipd_RAD2              : VitalDelayType01      := (0.0 ns, 0.0 ns);
        tipd_RAD1              : VitalDelayType01      := (0.0 ns, 0.0 ns);
        tipd_RAD0              : VitalDelayType01      := (0.0 ns, 0.0 ns);
tpd_WRAD4_WRDATA0         :VitalDelayType01Z := (2.0 ns,2.0 ns,2.0 ns,2.0 ns,2.0 ns,2.0 ns);
tpd_WRAD3_WRDATA0         :VitalDelayType01Z := (2.0 ns,2.0 ns,2.0 ns,2.0 ns,2.0 ns,2.0 ns);
tpd_WRAD2_WRDATA0         :VitalDelayType01Z := (2.0 ns,2.0 ns,2.0 ns,2.0 ns,2.0 ns,2.0 ns);
tpd_WRAD1_WRDATA0         :VitalDelayType01Z := (2.0 ns,2.0 ns,2.0 ns,2.0 ns,2.0 ns,2.0 ns);
tpd_WRAD0_WRDATA0         :VitalDelayType01Z := (2.0 ns,2.0 ns,2.0 ns,2.0 ns,2.0 ns,2.0 ns);
tpd_WRAD4_WRDATA1         :VitalDelayType01Z := (2.0 ns,2.0 ns,2.0 ns,2.0 ns,2.0 ns,2.0 ns);
tpd_WRAD3_WRDATA1         :VitalDelayType01Z := (2.0 ns,2.0 ns,2.0 ns,2.0 ns,2.0 ns,2.0 ns);
tpd_WRAD2_WRDATA1         :VitalDelayType01Z := (2.0 ns,2.0 ns,2.0 ns,2.0 ns,2.0 ns,2.0 ns);
tpd_WRAD1_WRDATA1         :VitalDelayType01Z := (2.0 ns,2.0 ns,2.0 ns,2.0 ns,2.0 ns,2.0 ns);
tpd_WRAD0_WRDATA1         :VitalDelayType01Z := (2.0 ns,2.0 ns,2.0 ns,2.0 ns,2.0 ns,2.0 ns);
tpd_WRAD4_WRDATA2         :VitalDelayType01Z := (2.0 ns,2.0 ns,2.0 ns,2.0 ns,2.0 ns,2.0 ns);
tpd_WRAD3_WRDATA2         :VitalDelayType01Z := (2.0 ns,2.0 ns,2.0 ns,2.0 ns,2.0 ns,2.0 ns);
tpd_WRAD2_WRDATA2         :VitalDelayType01Z := (2.0 ns,2.0 ns,2.0 ns,2.0 ns,2.0 ns,2.0 ns);
tpd_WRAD1_WRDATA2         :VitalDelayType01Z := (2.0 ns,2.0 ns,2.0 ns,2.0 ns,2.0 ns,2.0 ns);
tpd_WRAD0_WRDATA2         :VitalDelayType01Z := (2.0 ns,2.0 ns,2.0 ns,2.0 ns,2.0 ns,2.0 ns);
tpd_WRAD4_WRDATA3         :VitalDelayType01Z := (2.0 ns,2.0 ns,2.0 ns,2.0 ns,2.0 ns,2.0 ns);
tpd_WRAD3_WRDATA3         :VitalDelayType01Z := (2.0 ns,2.0 ns,2.0 ns,2.0 ns,2.0 ns,2.0 ns);
tpd_WRAD2_WRDATA3         :VitalDelayType01Z := (2.0 ns,2.0 ns,2.0 ns,2.0 ns,2.0 ns,2.0 ns);
tpd_WRAD1_WRDATA3         :VitalDelayType01Z := (2.0 ns,2.0 ns,2.0 ns,2.0 ns,2.0 ns,2.0 ns);
tpd_WRAD0_WRDATA3         :VitalDelayType01Z := (2.0 ns,2.0 ns,2.0 ns,2.0 ns,2.0 ns,2.0 ns);
tpd_OE_WRDATA0         :VitalDelayType01Z := (2.0 ns,2.0 ns,2.0 ns,2.0 ns,2.0 ns,2.0 ns);
tpd_OE_WRDATA1         :VitalDelayType01Z := (2.0 ns,2.0 ns,2.0 ns,2.0 ns,2.0 ns,2.0 ns);
tpd_OE_WRDATA2         :VitalDelayType01Z := (2.0 ns,2.0 ns,2.0 ns,2.0 ns,2.0 ns,2.0 ns);
tpd_OE_WRDATA3         :VitalDelayType01Z := (2.0 ns,2.0 ns,2.0 ns,2.0 ns,2.0 ns,2.0 ns);
tpd_ADRCLK_RDATA0         :VitalDelayType01 := (2.0 ns,2.0 ns);
tpd_ADRCLK_RDATA1         :VitalDelayType01 := (2.0 ns,2.0 ns);
tpd_ADRCLK_RDATA2         :VitalDelayType01 := (2.0 ns,2.0 ns);
tpd_ADRCLK_RDATA3         :VitalDelayType01 := (2.0 ns,2.0 ns);
tsetup_WRDATA3_WRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
thold_WRDATA3_WRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
tsetup_WRDATA2_WRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
thold_WRDATA2_WRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
tsetup_WRDATA1_WRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
thold_WRDATA1_WRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
tsetup_WRDATA0_WRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
thold_WRDATA0_WRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
tsetup_WRAD4_WRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
thold_WRAD4_WRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
tsetup_WRAD3_WRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
thold_WRAD3_WRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
tsetup_WRAD2_WRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
thold_WRAD2_WRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
tsetup_WRAD1_WRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
thold_WRAD1_WRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
tsetup_WRAD0_WRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
thold_WRAD0_WRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
tpw_WRCLK_posedge        :VitalDelayType := 1.0 ns;
tpw_ADRCLK_posedge        :VitalDelayType := 1.0 ns;
tsetup_WEN_ADRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
thold_WEN_ADRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
tsetup_RAD4_ADRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
thold_RAD4_ADRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
tsetup_RAD3_ADRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
thold_RAD3_ADRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
tsetup_RAD2_ADRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
thold_RAD2_ADRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
tsetup_RAD1_ADRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
thold_RAD1_ADRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
tsetup_RAD0_ADRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
thold_RAD0_ADRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
 
 
	TimingChecksOn : BOOLEAN := TRUE; 
	InstancePath : STRING := "*" 
            ); 
  PORT	( 
	WEN		: IN	std_logic ; 
	REN		: IN	std_logic ; 
	WRCLK		: IN	std_logic ; 
	ADRCLK		: IN	std_logic ; 
	OE		: IN	std_logic ; 
        WRDATA3         : INOUT std_logic := 'Z';
        WRDATA2         : INOUT std_logic := 'Z';
        WRDATA1         : INOUT std_logic := 'Z';
        WRDATA0         : INOUT std_logic := 'Z';
        RDATA3          :OUT std_logic := 'Z';
        RDATA2          : OUT std_logic := 'Z';
        RDATA1          : OUT std_logic := 'Z';
        RDATA0          : OUT std_logic := 'Z';
        RAD4           : IN    std_logic;
        RAD3           : IN    std_logic;
        RAD2           : IN    std_logic;
        RAD1           : IN    std_logic;
        RAD0           : IN    std_logic;
        WRAD4           : IN    std_logic;
        WRAD3           : IN    std_logic;
        WRAD2           : IN    std_logic;
        WRAD1           : IN    std_logic;
        WRAD0           : IN    std_logic
	); 
 
 
   ATTRIBUTE VITAL_LEVEL0 OF RB_DAR : ENTITY IS TRUE; 
 
END RB_DAR; 
 
----------------------------------------------------------------------- 
-- ARCHITECTURE declaration 
----------------------------------------------------------------------- 
ARCHITECTURE VITAL_VF OF RB_DAR IS 
 
    ATTRIBUTE VITAL_LEVEL1 OF VITAL_VF : ARCHITECTURE IS FALSE; 
 
	SIGNAL WEN_ipd		: std_logic := 'X'; 
	SIGNAL REN_ipd		: std_logic := 'X'; 
	SIGNAL WRCLK_ipd		: std_logic := '0'; 
	SIGNAL ADRCLK_ipd		: std_logic := '0'; 
	SIGNAL WR_CLK		: std_logic := '0'; 
	SIGNAL ADR_CLK		: std_logic := '0'; 
	SIGNAL OE_ipd	: std_logic := 'X'; 
	SIGNAL DIN		: std_logic_vector(3 DOWNTO 0); 
	SIGNAL RD_ADD		: std_logic_vector(4 DOWNTO 0); 
	SIGNAL r_add		: std_logic_vector(4 DOWNTO 0); 
	SIGNAL RD_ADD_W		: std_logic_vector(4 DOWNTO 0); 
	SIGNAL r_add_w		: std_logic_vector(4 DOWNTO 0); 
	SIGNAL WR_ADD		: std_logic_vector(4 DOWNTO 0); 
        SIGNAL WRDATA3_ipd      : std_logic := 'Z';
        SIGNAL WRDATA2_ipd      : std_logic := 'Z';
        SIGNAL WRDATA1_ipd      : std_logic := 'Z';
        SIGNAL WRDATA0_ipd      : std_logic := 'Z';
        SIGNAL WRAD4_ipd                : std_logic := '0';
        SIGNAL WRAD3_ipd                : std_logic := '0';
        SIGNAL WRAD2_ipd                : std_logic := '0';
        SIGNAL WRAD1_ipd                : std_logic := '0';
        SIGNAL WRAD0_ipd                : std_logic := '0';
        SIGNAL RAD4_ipd                : std_logic := '0';
        SIGNAL RAD3_ipd                : std_logic := '0';
        SIGNAL RAD2_ipd                : std_logic := '0';
        SIGNAL RAD1_ipd                : std_logic := '0';
        SIGNAL RAD0_ipd                : std_logic := '0';
	SIGNAL write_add	: std_logic_vector(4 DOWNTO 0); 
	SIGNAL data_out		: std_logic_vector(3 DOWNTO 0) := x_data; 
	SIGNAL data_out_w		: std_logic_vector(3 DOWNTO 0) := z_data; 
	SIGNAL output_delay	: time		:= 0 ns; 
	SIGNAL output_delay_w	: time		:= 0 ns; 
	SIGNAL memory_array	: memory_array_typ; 
 
BEGIN 
    
  --------------------------------------------------------------------- 
  -- INPUT PATH DELAYs 
  --------------------------------------------------------------------- 
  WIREDELAY : BLOCK 
  BEGIN 
	VitalWireDelay (WEN_ipd,		WEN,		tipd_WEN); 
	VitalWireDelay (REN_ipd,		REN,		tipd_REN); 
	VitalWireDelay (WRCLK_ipd,		WRCLK,		tipd_WRCLK); 
	VitalWireDelay (ADRCLK_ipd,		ADRCLK,		tipd_ADRCLK); 
	VitalWireDelay (OE_ipd,		OE,		tipd_OE); 
        VitalWireDelay (WRDATA0_ipd,    WRDATA0,        tipd_WRDATA0);
        VitalWireDelay (WRDATA1_ipd,    WRDATA1,        tipd_WRDATA1);
        VitalWireDelay (WRDATA2_ipd,    WRDATA2,        tipd_WRDATA2);
        VitalWireDelay (WRDATA3_ipd,    WRDATA3,        tipd_WRDATA3);
        VitalWireDelay (RAD0_ipd,              RAD0,          tipd_RAD0);
        VitalWireDelay (RAD1_ipd,              RAD1,          tipd_RAD1);
        VitalWireDelay (RAD2_ipd,              RAD2,          tipd_RAD2);
        VitalWireDelay (RAD3_ipd,              RAD3,          tipd_RAD3);
        VitalWireDelay (RAD4_ipd,              RAD4,          tipd_RAD4);
        VitalWireDelay (WRAD0_ipd,              WRAD0,          tipd_WRAD0);
        VitalWireDelay (WRAD1_ipd,              WRAD1,          tipd_WRAD1);
        VitalWireDelay (WRAD2_ipd,              WRAD2,          tipd_WRAD2);
        VitalWireDelay (WRAD3_ipd,              WRAD3,          tipd_WRAD3);
        VitalWireDelay (WRAD4_ipd,              WRAD4,          tipd_WRAD4); 
  END BLOCK; 
 
  --------------------------------------------------------------------- 
  -- Behavior Section 
  --------------------------------------------------------------------- 
 
  --------------------------------------------------------------------- 
  -- Wrapper Section 
  --------------------------------------------------------------------- 
 
   wrapper_latch_add_w : process(ADRCLK_ipd)
   
   begin
      if (ADRCLK_ipd = '1') then
           r_add_w(4) <= WRAD4_ipd;
           r_add_w(3) <= WRAD3_ipd;
           r_add_w(2) <= WRAD2_ipd;
           r_add_w(1) <= WRAD1_ipd;
           r_add_w(0) <= WRAD0_ipd;
      end if;

   end process;

  wrapper_latch_add : process(ADRCLK_ipd)
 
   begin
       if (ADRCLK_ipd = '1') then
           r_add(4) <= RAD4_ipd;
           r_add(3) <= RAD3_ipd;
           r_add(2) <= RAD2_ipd;
           r_add(1) <= RAD1_ipd;
           r_add(0) <= RAD0_ipd;
       end if;
  end process;
  
   wrapper_read_add : process(r_add, r_add_w) 
 
   begin 
	RD_ADD <= r_add; 
 
	RD_ADD_W <= r_add_w; 
   end process; 
 
   wrapper_write_add : process(WEN_ipd, WRAD4_ipd, WRAD3_ipd, WRAD2_ipd, WRAD1_ipd, WRAD0_ipd) 
 
   begin 
    if (WEN_ipd = '1') then 
        WR_ADD(4) <= WRAD4_ipd;
        WR_ADD(3) <= WRAD3_ipd;
        WR_ADD(2) <= WRAD2_ipd;
        WR_ADD(1) <= WRAD1_ipd;
        WR_ADD(0) <= WRAD0_ipd;
    else 
	WR_ADD <= x_add; 
    end if; 
 
   end process; 
 
   wrapper_write_clk : process(WEN_ipd, WRCLK_ipd) 
 
   begin 
    if (WEN_ipd = '1') then 
	WR_CLK <= WRCLK_ipd; 
    else 
	WR_CLK <= '0'; 
    end if; 
 
   end process; 

   wrapper_addr_clk : process(ADRCLK_ipd,WEN_ipd) 
 
   begin 
      if (WEN_ipd = '0') then
	ADR_CLK <= ADRCLK_ipd; 
      else
        ADR_CLK <= '0';
      end if;
    end process; 
 
   process(WR_CLK) 
 
    begin 
      if WR_CLK = '1' then 
        write_add(4) <= WRAD4_ipd;
        write_add(3) <= WRAD3_ipd;
        write_add(2) <= WRAD2_ipd;
        write_add(1) <= WRAD1_ipd;
        write_add(0) <= WRAD0_ipd;
      end if; 
 
   end process; 
 
   wrapper_write_data : process(WEN_ipd, WRDATA3_ipd, WRDATA2_ipd, WRDATA1_ipd, WRDATA0_ipd) 
 
   begin 
    if (WEN_ipd = '1') then 
        DIN(3) <= WRDATA3_ipd;
        DIN(2) <= WRDATA2_ipd;
        DIN(1) <= WRDATA1_ipd;
        DIN(0) <= WRDATA0_ipd;
    else 
	DIN <= x_data; 
    end if; 
 
   end process; 
 
 
  VITALBehavior : PROCESS ( WEN_ipd, REN_ipd, WR_CLK, ADRCLK, ADR_CLK,  DIN, RD_ADD_W, RD_ADD, WR_ADD, RAD4_ipd, RAD3_ipd, RAD2_ipd, RAD1_ipd, RAD0_ipd ) 
 
 
   -- Temporary variables 
   VARIABLE tempaddr 		: integer := 0; 
   VARIABLE rd_address 		: integer := 0; 
   VARIABLE rd_address_w 	: integer := 0; 
   VARIABLE rd_viol_flag 	: X01 := '0'; 
   VARIABLE rd_viol_flag_w 	: X01 := '0'; 
 
   -- Timing Check results 
   VARIABLE Pviol_WRCLK			: std_logic := '0'; 
   VARIABLE PeriodData_WRCLK		: VitalPeriodDataType := VitalPeriodDataInit; 
   VARIABLE Pviol_ADRCLK			: std_logic := '0'; 
   VARIABLE PeriodData_ADRCLK		: VitalPeriodDataType := VitalPeriodDataInit; 
   VARIABLE Tviol_WR_ADD_stp_hld_0	: std_logic := '0'; 
   VARIABLE TimingData_WR_ADD_stp_hld_0	: VitalTimingDataType := VitalTimingDataInit; 
   VARIABLE Tviol_WR_ADD_stp_hld_1	: std_logic := '0'; 
   VARIABLE TimingData_WR_ADD_stp_hld_1	: VitalTimingDataType := VitalTimingDataInit; 
   VARIABLE Tviol_WR_ADD_stp_hld_2	: std_logic := '0'; 
   VARIABLE TimingData_WR_ADD_stp_hld_2	: VitalTimingDataType := VitalTimingDataInit; 
   VARIABLE Tviol_WR_ADD_stp_hld_3	: std_logic := '0'; 
   VARIABLE TimingData_WR_ADD_stp_hld_3	: VitalTimingDataType := VitalTimingDataInit; 
   VARIABLE Tviol_WR_ADD_stp_hld_4	: std_logic := '0'; 
   VARIABLE TimingData_WR_ADD_stp_hld_4	: VitalTimingDataType := VitalTimingDataInit; 
   VARIABLE Tviol_WR_DATA_stp_0		: std_logic := '0'; 
   VARIABLE TimingData_WR_DATA_stp_0	: VitalTimingDataType := VitalTimingDataInit; 
   VARIABLE Tviol_WR_DATA_stp_1		: std_logic := '0'; 
   VARIABLE TimingData_WR_DATA_stp_1	: VitalTimingDataType := VitalTimingDataInit; 
   VARIABLE Tviol_WR_DATA_stp_2		: std_logic := '0'; 
   VARIABLE TimingData_WR_DATA_stp_2	: VitalTimingDataType := VitalTimingDataInit; 
   VARIABLE Tviol_WR_DATA_stp_3		: std_logic := '0'; 
   VARIABLE TimingData_WR_DATA_stp_3	: VitalTimingDataType := VitalTimingDataInit; 
   VARIABLE Tviol_WR_DATA_hld_0		: std_logic := '0'; 
   VARIABLE TimingData_WR_DATA_hld_0	: VitalTimingDataType := VitalTimingDataInit; 
   VARIABLE Tviol_WR_DATA_hld_1		: std_logic := '0'; 
   VARIABLE TimingData_WR_DATA_hld_1	: VitalTimingDataType := VitalTimingDataInit; 
   VARIABLE Tviol_WR_DATA_hld_2		: std_logic := '0'; 
   VARIABLE TimingData_WR_DATA_hld_2	: VitalTimingDataType := VitalTimingDataInit; 
   VARIABLE Tviol_WR_DATA_hld_3		: std_logic := '0'; 
   VARIABLE TimingData_WR_DATA_hld_3	: VitalTimingDataType := VitalTimingDataInit; 
   VARIABLE Tviol_RD_ADD_stp_hld_0		: std_logic := '0'; 
   VARIABLE TimingData_RD_ADD_stp_hld_0	: VitalTimingDataType := VitalTimingDataInit; 
   VARIABLE Tviol_RD_ADD_stp_hld_1		: std_logic := '0'; 
   VARIABLE TimingData_RD_ADD_stp_hld_1	: VitalTimingDataType := VitalTimingDataInit; 
   VARIABLE Tviol_RD_ADD_stp_hld_2		: std_logic := '0'; 
   VARIABLE TimingData_RD_ADD_stp_hld_2	: VitalTimingDataType := VitalTimingDataInit; 
   VARIABLE Tviol_RD_ADD_stp_hld_3		: std_logic := '0'; 
   VARIABLE TimingData_RD_ADD_stp_hld_3	: VitalTimingDataType := VitalTimingDataInit; 
   VARIABLE Tviol_RD_ADD_stp_hld_4		: std_logic := '0'; 
   VARIABLE TimingData_RD_ADD_stp_hld_4	: VitalTimingDataType := VitalTimingDataInit; 
   VARIABLE Tviol_WEN_hld		: std_logic := '0'; 
   VARIABLE TimingData_WEN_hld		: VitalTimingDataType := VitalTimingDataInit; 
 
 
 
 BEGIN 
    ------------------------------------------------------------------- 
    -- Timing Check Section 
    ------------------------------------------------------------------- 
    IF (TimingChecksOn) THEN 
 
	VitalPeriodPulseCheck  (Pviol_WRCLK, 
				PeriodData_WRCLK, 
				WR_CLK, "WRCLK", 
				0.0 ns, 
				0.0 ns, 
				tpw_WRCLK_posedge, 
				0.0 ns, 
				True,
				InstancePath & "/RB_DAR", 
				TRUE, 
				TRUE, 
				WARNING ); 

	VitalPeriodPulseCheck  (Pviol_ADRCLK, 
				PeriodData_ADRCLK, 
				ADR_CLK, "ADRCLK", 
				0.0 ns, 
				0.0 ns, 
				tpw_ADRCLK_posedge, 
				0.0 ns, 
				True,
				InstancePath & "/RB_DAR", 
				TRUE, 
				TRUE, 
				WARNING ); 
 
        VitalSetupHoldCheck    (Tviol_WR_ADD_stp_hld_0,
                                TimingData_WR_ADD_stp_hld_0,
                                WR_ADD(0), "WRAD0",
                                0.0 ns,
                                WR_CLK, "WRCLK",
                                0.0 ns,
                                tsetup_WRAD0_WRCLK_noedge_posedge, tsetup_WRAD0_WRCLK_noedge_posedge,
                                thold_WRAD0_WRCLK_noedge_posedge, thold_WRAD0_WRCLK_noedge_posedge,
                                WEN_ipd = '1',
                                '/',
                                InstancePath & "/RB_DAR",
                                TRUE,
                                TRUE,
                                WARNING );

        VitalSetupHoldCheck    (Tviol_WR_ADD_stp_hld_1,
                                TimingData_WR_ADD_stp_hld_1,
                                WR_ADD(1), "WRAD1",
                                0.0 ns,
                                WR_CLK, "WRCLK",
                                0.0 ns,
                                tsetup_WRAD1_WRCLK_noedge_posedge, tsetup_WRAD1_WRCLK_noedge_posedge,
                                thold_WRAD1_WRCLK_noedge_posedge, thold_WRAD1_WRCLK_noedge_posedge,
                                WEN_ipd = '1',
                                '/',
                                InstancePath & "/RB_DAR",
                                TRUE,
                                TRUE,
                                WARNING );

        VitalSetupHoldCheck    (Tviol_WR_ADD_stp_hld_2,
                                TimingData_WR_ADD_stp_hld_2,
                                WR_ADD(2), "WRAD2",
                                0.0 ns,
                                WR_CLK, "WRCLK",
                                0.0 ns,
                                tsetup_WRAD2_WRCLK_noedge_posedge, tsetup_WRAD2_WRCLK_noedge_posedge,
                                thold_WRAD2_WRCLK_noedge_posedge, thold_WRAD2_WRCLK_noedge_posedge,
                                WEN_ipd = '1',
                                '/',
                                InstancePath & "/RB_DAR",
                                TRUE,
                                TRUE,
                                WARNING );
       VitalSetupHoldCheck    (Tviol_WR_ADD_stp_hld_3,
                                TimingData_WR_ADD_stp_hld_3,
                                WR_ADD(3), "WRAD3",
                                0.0 ns,
                                WR_CLK, "WRCLK",
                                0.0 ns,
                                tsetup_WRAD3_WRCLK_noedge_posedge, tsetup_WRAD3_WRCLK_noedge_posedge,
                                thold_WRAD3_WRCLK_noedge_posedge, thold_WRAD3_WRCLK_noedge_posedge,
                                WEN_ipd = '1',
                                '/',
                                InstancePath & "/RB_DAR",
                                TRUE,
                                TRUE,
                                WARNING );
  VitalSetupHoldCheck    (Tviol_WR_ADD_stp_hld_4,
                                TimingData_WR_ADD_stp_hld_4,
                                WR_ADD(4), "WRAD4",
                                0.0 ns,
                                WR_CLK, "WRCLK",
                                0.0 ns,
                                tsetup_WRAD4_WRCLK_noedge_posedge, tsetup_WRAD4_WRCLK_noedge_posedge,
                                thold_WRAD4_WRCLK_noedge_posedge, thold_WRAD4_WRCLK_noedge_posedge,
                                WEN_ipd = '1',
                                '/',
                                InstancePath & "/RB_DAR",
                                TRUE,
                                TRUE,
                                WARNING );

        VitalSetupHoldCheck    (Tviol_WR_DATA_stp_0,
                                TimingData_WR_DATA_stp_0,
                                DIN(0), "WRDATA0",
                                0.0 ns,
                                WR_CLK, "WRCLK",
                                0.0 ns,
                                tsetup_WRDATA0_WRCLK_noedge_posedge, tsetup_WRDATA0_WRCLK_noedge_posedge,
                                0.0 ns, 0.0 ns,
                                WEN_ipd = '1',
                                '/',
                                InstancePath & "/RB_DAR",
                                TRUE,
                                TRUE,
                                WARNING );

        VitalSetupHoldCheck    (Tviol_WR_DATA_stp_1,
                                TimingData_WR_DATA_stp_1,
                                DIN(1), "WRDATA1",
                                0.0 ns,
                                WR_CLK, "WRCLK",
                                0.0 ns,
                                tsetup_WRDATA1_WRCLK_noedge_posedge, tsetup_WRDATA1_WRCLK_noedge_posedge,
                                0.0 ns, 0.0 ns,
                                WEN_ipd = '1',
                                '/',
                                InstancePath & "/RB_DAR",
                                TRUE,
                                TRUE,
                                WARNING );

        VitalSetupHoldCheck    (Tviol_WR_DATA_stp_2,
                                TimingData_WR_DATA_stp_2,
                                DIN(2), "WRDATA2",
                                0.0 ns,
                                WR_CLK, "WRCLK",
                                0.0 ns,
                                tsetup_WRDATA2_WRCLK_noedge_posedge, tsetup_WRDATA2_WRCLK_noedge_posedge,
                                0.0 ns, 0.0 ns,
                                WEN_ipd = '1',
                                '/',
                                InstancePath & "/RB_DAR",
                                TRUE,
                                TRUE,
                                WARNING );
        VitalSetupHoldCheck    (Tviol_WR_DATA_stp_3,
                                TimingData_WR_DATA_stp_3,
                                DIN(3), "WRDATA3",
                                0.0 ns,
                                WR_CLK, "WRCLK",
                                0.0 ns,
                                tsetup_WRDATA3_WRCLK_noedge_posedge, tsetup_WRDATA3_WRCLK_noedge_posedge,
                                0.0 ns, 0.0 ns,
                                WEN_ipd = '1',
                                '/',
                                InstancePath & "/RB_DAR",
                                TRUE,
                                TRUE,
                                WARNING );

        VitalSetupHoldCheck    (Tviol_WR_DATA_hld_0,
                                TimingData_WR_DATA_hld_0,
                                DIN(0), "WRDATA0",
                                0.0 ns,
                                WR_CLK, "WRCLK",
                                0.0 ns,
                                0.0 ns, 0.0 ns,
                                thold_WRDATA0_WRCLK_noedge_posedge, thold_WRDATA0_WRCLK_noedge_posedge,
                                WEN_ipd = '1',
                                '/',
                                InstancePath & "/RB_DAR",
                                TRUE,
                                TRUE,
                                WARNING );

        VitalSetupHoldCheck    (Tviol_WR_DATA_hld_1,
                                TimingData_WR_DATA_hld_1,
                                DIN(1), "WRDATA1",
                                0.0 ns,
                                WR_CLK, "WRCLK",
                                0.0 ns,
                                0.0 ns, 0.0 ns,
                                thold_WRDATA1_WRCLK_noedge_posedge, thold_WRDATA1_WRCLK_noedge_posedge,
                                WEN_ipd = '1',
                                '/',
                                InstancePath & "/RB_DAR",
                                TRUE,
                                TRUE,
                                WARNING );

        VitalSetupHoldCheck    (Tviol_WR_DATA_hld_2,
                                TimingData_WR_DATA_hld_2,
                                DIN(2), "WRDATA2",
                                0.0 ns,
                                WR_CLK, "WRCLK",
                                0.0 ns,
                                0.0 ns, 0.0 ns,
                                thold_WRDATA2_WRCLK_noedge_posedge, thold_WRDATA2_WRCLK_noedge_posedge,
                                WEN_ipd = '1',
                                '/',
                                InstancePath & "/RB_DAR",
                                TRUE,
                                TRUE,
                                WARNING );
        VitalSetupHoldCheck    (Tviol_WR_DATA_hld_3,
                                TimingData_WR_DATA_hld_3,
                                DIN(3), "WRDATA3",
                                0.0 ns,
                                WR_CLK, "WRCLK",
                                0.0 ns,
                                0.0 ns, 0.0 ns,
                                thold_WRDATA3_WRCLK_noedge_posedge, thold_WRDATA3_WRCLK_noedge_posedge,
                                WEN_ipd = '1',
                                '/',
                                InstancePath & "/RB_DAR",
                                TRUE,
                                TRUE,
                                WARNING );
        VitalSetupHoldCheck    (Tviol_RD_ADD_stp_hld_0,
                                TimingData_RD_ADD_stp_hld_0,
                                RAD0_ipd, "RAD0",
                                0.0 ns,
                                ADRCLK_ipd, "ADRCLK",
                                0.0 ns,
                                tsetup_RAD0_ADRCLK_noedge_posedge, tsetup_RAD0_ADRCLK_noedge_posedge,
                                thold_RAD0_ADRCLK_noedge_posedge, thold_RAD0_ADRCLK_noedge_posedge,
                                True,
                                '/',
                                InstancePath & "/RB_DAR",
                                TRUE,
                                TRUE,
                                WARNING );

        VitalSetupHoldCheck    (Tviol_RD_ADD_stp_hld_1,
                                TimingData_RD_ADD_stp_hld_1,
                                RAD1_ipd, "RAD1",
                                0.0 ns,
                                ADRCLK_ipd, "ADRCLK",
                                0.0 ns,
                                tsetup_RAD1_ADRCLK_noedge_posedge, tsetup_RAD1_ADRCLK_noedge_posedge,
                                thold_RAD1_ADRCLK_noedge_posedge, thold_RAD1_ADRCLK_noedge_posedge,
                                True,
                                '/',
                                InstancePath & "/RB_DAR",
                                TRUE,
                                TRUE,
                                WARNING );

        VitalSetupHoldCheck    (Tviol_RD_ADD_stp_hld_2,
                                TimingData_RD_ADD_stp_hld_2,
                                RAD2_ipd, "RAD2",
                                0.0 ns,
                                ADRCLK_ipd, "ADRCLK",
                                0.0 ns,
                                tsetup_RAD2_ADRCLK_noedge_posedge, tsetup_RAD2_ADRCLK_noedge_posedge,
                                thold_RAD2_ADRCLK_noedge_posedge, thold_RAD2_ADRCLK_noedge_posedge,
                                True,
                                '/',
                                InstancePath & "/RB_DAR",
                                TRUE,
                                TRUE,
                                WARNING );

        VitalSetupHoldCheck    (Tviol_RD_ADD_stp_hld_3,
                                TimingData_RD_ADD_stp_hld_3,
                                RAD3_ipd, "RAD3",
                                0.0 ns,
                                ADRCLK_ipd, "ADRCLK",
                                0.0 ns,
                                tsetup_RAD3_ADRCLK_noedge_posedge, tsetup_RAD3_ADRCLK_noedge_posedge,
                                thold_RAD3_ADRCLK_noedge_posedge, thold_RAD3_ADRCLK_noedge_posedge,
                                True,
                                '/',
                                InstancePath & "/RB_DAR",
                                TRUE,
                                TRUE,
                                WARNING );
        VitalSetupHoldCheck    (Tviol_RD_ADD_stp_hld_4,
                                TimingData_RD_ADD_stp_hld_4,
                                RAD4_ipd, "RAD4",
                                0.0 ns,
                                ADRCLK_ipd, "ADRCLK",
                                0.0 ns,
                                tsetup_RAD4_ADRCLK_noedge_posedge, tsetup_RAD4_ADRCLK_noedge_posedge,
                                thold_RAD4_ADRCLK_noedge_posedge, thold_RAD4_ADRCLK_noedge_posedge,
                                True,
                                '/',
                                InstancePath & "/RB_DAR",
                                TRUE,
                                TRUE,
                                WARNING );

	VitalSetupHoldCheck    (Tviol_WEN_hld, 
				TimingData_WEN_hld, 
				WEN_ipd, "WEN", 
				0.0 ns, 
				ADR_CLK, "ADRCLK", 
				0.0 ns, 
				tsetup_WEN_ADRCLK_noedge_posedge, tsetup_WEN_ADRCLK_noedge_posedge,
				thold_WEN_ADRCLK_noedge_posedge, thold_WEN_ADRCLK_noedge_posedge,
				True, 
				'/', 
				InstancePath & "/RB_DAR", 
				TRUE, 
				TRUE, 
				WARNING ); 
 
    END IF; -- Timing Check Section 

 
 rd_viol_flag :=  (Tviol_RD_ADD_stp_hld_0 or Tviol_RD_ADD_stp_hld_1 or Tviol_RD_ADD_stp_hld_2 or Tviol_RD_ADD_stp_hld_3 or Tviol_RD_ADD_stp_hld_4 or Pviol_ADRCLK); 

 
 
 
    ------------------------------------------------------------------- 
    -- Functionality Section 
    ------------------------------------------------------------------- 
 
-- WRITE ADDRESS GOES XX 
 
    if ( WR_CLK'EVENT and WR_CLK = '1' and vecX(WR_ADD)) then 
 
        assert false 
        report "Illegal Address Input: Undefined  Address at the Read_Write Port." 
        severity note ; 
        memory_array <= (others => x_data); 
 
    end if; 
 
-- ADDRESS HOLD AND SETUP VIOLATION EFFECT 
 
    if( Tviol_WR_ADD_stp_hld_0 = 'X' or Tviol_WR_ADD_stp_hld_1 = 'X' or Tviol_WR_ADD_stp_hld_2 = 'X' or Tviol_WR_ADD_stp_hld_3 = 'X' or Tviol_WR_ADD_stp_hld_4 = 'X' ) then 
 
        memory_array <= (others => x_data); 
 
    else 
 
-- DATA SETUP AND HOLD VIOLATION EFFECT 
 
    if( Pviol_WRCLK = 'X' or Tviol_WR_DATA_hld_0 = 'X' or Tviol_WR_DATA_hld_1 = 'X' or Tviol_WR_DATA_hld_2 = 'X' or Tviol_WR_DATA_hld_3 = 'X' or Tviol_WEN_hld = 'X') then 
	tempaddr := vec2int(write_add); 
	memory_array(tempaddr) <= x_data; 
    end if; 
 
    if( Tviol_WR_DATA_stp_0 = 'X' or Tviol_WR_DATA_stp_1 = 'X' or Tviol_WR_DATA_stp_2 = 'X' or Tviol_WR_DATA_stp_3 = 'X') then 
	tempaddr := vec2int(WR_ADD); 
	memory_array(tempaddr) <= x_data; 
    end if; 
 
    end if; 
 
-- VALID MEMORY WRITE 
 
    if ( WR_CLK'EVENT and WR_CLK = '1' and not(vecX(WR_ADD)) and not(Tviol_WR_ADD_stp_hld_0 = 'X' or Tviol_WR_ADD_stp_hld_1 = 'X' or Tviol_WR_ADD_stp_hld_2 = 'X' or Tviol_WR_ADD_stp_hld_3 = 'X' or Tviol_WR_ADD_stp_hld_4 = 'X') and not( Pviol_WRCLK = 'X' or Tviol_WR_DATA_hld_0 = 'X' or Tviol_WR_DATA_hld_1 = 'X' or Tviol_WR_DATA_hld_2 = 'X' or Tviol_WR_DATA_hld_3 = 'X' or Tviol_WEN_hld = 'X') and not( Tviol_WR_DATA_stp_0 = 'X' or Tviol_WR_DATA_stp_1 = 'X' or Tviol_WR_DATA_stp_2 = 'X' or Tviol_WR_DATA_stp_3 = 'X')) then 
	tempaddr := vec2int(WR_ADD); 
	memory_array(tempaddr) <= DIN; 
    end if; 
 
    if WR_CLK'EVENT and WR_CLK /= WRCLK_ipd and WR_CLK'LAST_VALUE = '1' then 
	memory_array(tempaddr) <= x_data; 
    end if; 
 
 
-- READ CYCLE VIOLATION EFFECT 
 
    if( rd_viol_flag = 'X' or (RD_ADD'EVENT and REN_ipd = '1' and vecX(RD_ADD))) then 
	data_out <= x_data; 
    elsif 
 
-- VALID MEMORY READ 
 
     (RD_ADD'EVENT and REN_ipd = '1' and not(rd_viol_flag = 'X') and not (vecX(RD_ADD))) then 
	rd_address := vec2int(RD_ADD); 
	data_out <= TRANSPORT memory_array(rd_address); 
    end if; 
 
 
    if((RD_ADD_W'EVENT and REN_ipd = '1' and OE_ipd = '1' and vecX(RD_ADD_W))) then 
	data_out_w <= x_data; 
    elsif 
 
-- VALID MEMORY READ 
 
     (RD_ADD_W'EVENT  and REN_ipd = '1' and OE_ipd = '1' and WEN_ipd = '0' and not (vecX(RD_ADD_W))) then 
	rd_address_w := vec2int(RD_ADD_W); 
	data_out_w <= TRANSPORT memory_array(rd_address_w); 
    end if; 
 
  END PROCESS; 
 
    ------------------------------------------------------------------------------- 
    -- Temporary output signal should get assigned to the output signal. 
    ------------------------------------------------------------------------------- 
 
 
   PROCESS(data_out, data_out_w, REN_ipd, OE_ipd, ADRCLK_ipd, WRAD4_ipd, WRAD3_ipd, WRAD2_ipd, WRAD1_ipd, WRAD0_ipd)

   VARIABLE GLITCH_DATA : VitalGlitchDataType;
   VARIABLE GLITCH : VitalGlitchDataType;
   VARIABLE con : std_logic ;--:= '0';
    VARIABLE WEN_inv : std_logic ;--:= '0';
    VARIABLE WRDATA3_1 : std_logic := 'Z';
    VARIABLE WRDATA2_1 : std_logic := 'Z';
    VARIABLE WRDATA1_1 : std_logic := 'Z';
    VARIABLE WRDATA0_1 : std_logic := 'Z';
    VARIABLE RDATA3_1 : std_logic := 'X';
    VARIABLE RDATA2_1 : std_logic := 'X';
    VARIABLE RDATA1_1 : std_logic := 'X';
    VARIABLE RDATA0_1 : std_logic := 'X';

   BEGIN
       WEN_inv := VitalINV(WEN_ipd);
       con := VitalAND3(OE_ipd,REN_ipd, WEN_inv);


      WRDATA3_1 := VITALBUFIF1(data_out_w(3),con);
      WRDATA2_1 := VITALBUFIF1(data_out_w(2),con);
      WRDATA1_1 := VITALBUFIF1(data_out_w(1),con);
      WRDATA0_1 := VITALBUFIF1(data_out_w(0),con);

      RDATA3_1 := VITALBUF(data_out(3));
      RDATA2_1 := VITALBUF(data_out(2));
      RDATA1_1 := VITALBUF(data_out(1));
      RDATA0_1 := VITALBUF(data_out(0));

     VitalPathDelay01 ( RDATA3, GLITCH, "RDATA3", RDATA3_1,
        Paths => (
        0 => ( ADRCLK_ipd'LAST_EVENT, tpd_ADRCLK_RDATA3, TRUE )),
        DefaultDelay=>VitalZeroDelay01,
        Mode=>VitalInertial,
        XON=>TRUE,
        MsgOn=>TRUE,
        MsgSeverity=>WARNING );

     VitalPathDelay01 ( RDATA2, GLITCH, "RDATA2", RDATA2_1,
        Paths => (
        0 => ( ADRCLK_ipd'LAST_EVENT, tpd_ADRCLK_RDATA2, TRUE )),
        DefaultDelay=>VitalZeroDelay01,
        Mode=>VitalInertial,
        XON=>TRUE,
        MsgOn=>TRUE,
        MsgSeverity=>WARNING );

     VitalPathDelay01 ( RDATA1, GLITCH, "RDATA1", RDATA1_1,
        Paths => (
        0 => ( ADRCLK_ipd'LAST_EVENT, tpd_ADRCLK_RDATA1, TRUE )),
        DefaultDelay=>VitalZeroDelay01,
        Mode=>VitalInertial,
        XON=>TRUE,
        MsgOn=>TRUE,
        MsgSeverity=>WARNING );

     VitalPathDelay01 ( RDATA0, GLITCH, "RDATA0", RDATA0_1,
        Paths => (
        0 => ( ADRCLK_ipd'LAST_EVENT, tpd_ADRCLK_RDATA0, TRUE )),
        DefaultDelay=>VitalZeroDelay01,
        Mode=>VitalInertial,
        XON=>TRUE,
        MsgOn=>TRUE,
        MsgSeverity=>WARNING );


      VitalPathDelay01Z ( WRDATA3, GLITCH_DATA, "WRDATA3", WRDATA3_1,
        Paths => (
        0 => ( WRAD4_ipd'LAST_EVENT, VitalExtendToFillDelay(tpd_WRAD4_WRDATA3), TRUE ),
        1 => ( WRAD3_ipd'LAST_EVENT, VitalExtendToFillDelay(tpd_WRAD3_WRDATA3), TRUE ),
        2 => ( WRAD2_ipd'LAST_EVENT, VitalExtendToFillDelay(tpd_WRAD2_WRDATA3), TRUE ),
        3 => ( WRAD1_ipd'LAST_EVENT, VitalExtendToFillDelay(tpd_WRAD1_WRDATA3), TRUE ),
        4 => ( WRAD0_ipd'LAST_EVENT, VitalExtendToFillDelay(tpd_WRAD0_WRDATA3), TRUE ),
        5 => ( OE_ipd'LAST_EVENT, VitalExtendToFillDelay(tpd_OE_WRDATA3), TRUE ) ),
        DefaultDelay=>VitalZeroDelay01Z,
        Mode=>VitalInertial,
        XON=>TRUE,
        MsgOn=>TRUE,
        MsgSeverity=>WARNING,
        OutputMap => "UX01ZWLH-");

      VitalPathDelay01Z ( WRDATA2, GLITCH_DATA, "WRDATA2", WRDATA2_1,
        Paths => (
        0 => ( WRAD4_ipd'LAST_EVENT, VitalExtendToFillDelay(tpd_WRAD4_WRDATA2), TRUE ),
        1 => ( WRAD3_ipd'LAST_EVENT, VitalExtendToFillDelay(tpd_WRAD3_WRDATA2), TRUE ),
        2 => ( WRAD2_ipd'LAST_EVENT, VitalExtendToFillDelay(tpd_WRAD2_WRDATA2), TRUE ),
        3 => ( WRAD1_ipd'LAST_EVENT, VitalExtendToFillDelay(tpd_WRAD1_WRDATA2), TRUE ),
        4 => ( WRAD0_ipd'LAST_EVENT, VitalExtendToFillDelay(tpd_WRAD0_WRDATA2), TRUE ),
        5 => ( OE_ipd'LAST_EVENT, VitalExtendToFillDelay(tpd_OE_WRDATA2), TRUE ) ),
        DefaultDelay=>VitalZeroDelay01Z,
        Mode=>VitalInertial,
        XON=>TRUE,
        MsgOn=>TRUE,
        MsgSeverity=>WARNING,
        OutputMap => "UX01ZWLH-");

      VitalPathDelay01Z ( WRDATA1, GLITCH_DATA, "WRDATA1", WRDATA1_1,
        Paths => (
        0 => ( WRAD4_ipd'LAST_EVENT, VitalExtendToFillDelay(tpd_WRAD4_WRDATA1), TRUE ),
        1 => ( WRAD3_ipd'LAST_EVENT, VitalExtendToFillDelay(tpd_WRAD3_WRDATA1), TRUE ),
        2 => ( WRAD2_ipd'LAST_EVENT, VitalExtendToFillDelay(tpd_WRAD2_WRDATA1), TRUE ),
        3 => ( WRAD1_ipd'LAST_EVENT, VitalExtendToFillDelay(tpd_WRAD1_WRDATA1), TRUE ),
        4 => ( WRAD0_ipd'LAST_EVENT, VitalExtendToFillDelay(tpd_WRAD0_WRDATA1), TRUE ),
        5 => ( OE_ipd'LAST_EVENT, VitalExtendToFillDelay(tpd_OE_WRDATA1), TRUE ) ),
        DefaultDelay=>VitalZeroDelay01Z,
        Mode=>VitalInertial,
        XON=>TRUE,
        MsgOn=>TRUE,
        MsgSeverity=>WARNING,
        OutputMap => "UX01ZWLH-");

       VitalPathDelay01Z ( WRDATA0, GLITCH_DATA, "WRDATA0", WRDATA0_1,
        Paths => (
        0 => ( WRAD4_ipd'LAST_EVENT, VitalExtendToFillDelay(tpd_WRAD4_WRDATA0), TRUE ),
        1 => ( WRAD3_ipd'LAST_EVENT, VitalExtendToFillDelay(tpd_WRAD3_WRDATA0), TRUE ),
        2 => ( WRAD2_ipd'LAST_EVENT, VitalExtendToFillDelay(tpd_WRAD2_WRDATA0), TRUE ),
        3 => ( WRAD1_ipd'LAST_EVENT, VitalExtendToFillDelay(tpd_WRAD1_WRDATA0), TRUE ),
        4 => ( WRAD0_ipd'LAST_EVENT, VitalExtendToFillDelay(tpd_WRAD0_WRDATA0), TRUE ),
        5 => ( OE_ipd'LAST_EVENT, VitalExtendToFillDelay(tpd_OE_WRDATA0), TRUE ) ),
        DefaultDelay=>VitalZeroDelay01Z,
        Mode=>VitalInertial,
        XON=>TRUE,
        MsgOn=>TRUE,
        MsgSeverity=>WARNING,
        OutputMap => "UX01ZWLH-");

END PROCESS;
 
 
END VITAL_VF; 
configuration CFG_RB_DAR_VITAL of RB_DAR is
        for VITAL_VF
        end for;
end CFG_RB_DAR_VITAL;
----------------------------------------------------------------------- 
 
-- VITAL model for RB_MAR 30.10 technology 
----------------------------------------------------------------------- 
 
LIBRARY IEEE; 
USE IEEE.std_logic_1164.ALL; 
USE IEEE.VITAL_timing.all; 
USE IEEE.std_logic_textio.all; 
USE IEEE.VITAL_primitives.all; 
LIBRARY std; 
USE std.textio.all; 
LIBRARY VF1; 
USE VF1.ALL; 
USE VF1.RAMPACK.ALL; 
 
----------------------------------------------------------------------- 
-- ENTITY declaration 
----------------------------------------------------------------------- 
 
ENTITY RB_MAR IS 
  GENERIC ( 
	tipd_WEN		: VitalDelayType01			:= (0.0 ns, 0.0 ns); 
	tipd_WRCLK		: VitalDelayType01			:= (0.0 ns, 0.0 ns); 
	tipd_ADRCLK		: VitalDelayType01			:= (0.0 ns, 0.0 ns); 
	tipd_OE		: VitalDelayType01			:= (0.0 ns, 0.0 ns); 
        tipd_WRDATA3            : VitalDelayType01      := (0.0 ns, 0.0 ns);
        tipd_WRDATA2            : VitalDelayType01      := (0.0 ns, 0.0 ns);
        tipd_WRDATA1            : VitalDelayType01      := (0.0 ns, 0.0 ns);
        tipd_WRDATA0            : VitalDelayType01      := (0.0 ns, 0.0 ns);
        tipd_WRAD4              : VitalDelayType01      := (0.0 ns, 0.0 ns);
        tipd_WRAD3              : VitalDelayType01      := (0.0 ns, 0.0 ns);
        tipd_WRAD2              : VitalDelayType01      := (0.0 ns, 0.0 ns);
        tipd_WRAD1              : VitalDelayType01      := (0.0 ns, 0.0 ns);
        tipd_WRAD0              : VitalDelayType01      := (0.0 ns, 0.0 ns);
tpd_OE_WRDATA0         :VitalDelayType01Z := (2.0 ns,2.0 ns,2.0 ns,2.0 ns,2.0 ns,2.0 ns);
tpd_OE_WRDATA1         :VitalDelayType01Z := (2.0 ns,2.0 ns,2.0 ns,2.0 ns,2.0 ns,2.0 ns);
tpd_OE_WRDATA2         :VitalDelayType01Z := (2.0 ns,2.0 ns,2.0 ns,2.0 ns,2.0 ns,2.0 ns);
tpd_OE_WRDATA3         :VitalDelayType01Z := (2.0 ns,2.0 ns,2.0 ns,2.0 ns,2.0 ns,2.0 ns);
tpd_ADRCLK_WRDATA0         :VitalDelayType01Z := (2.0 ns,2.0 ns,2.0 ns,2.0 ns,2.0 ns,2.0 ns);
tpd_ADRCLK_WRDATA1         :VitalDelayType01Z := (2.0 ns,2.0 ns,2.0 ns,2.0 ns,2.0 ns,2.0 ns);
tpd_ADRCLK_WRDATA2         :VitalDelayType01Z := (2.0 ns,2.0 ns,2.0 ns,2.0 ns,2.0 ns,2.0 ns);
tpd_ADRCLK_WRDATA3         :VitalDelayType01Z := (2.0 ns,2.0 ns,2.0 ns,2.0 ns,2.0 ns,2.0 ns);
tsetup_WRDATA3_WRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
thold_WRDATA3_WRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
tsetup_WRDATA2_WRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
thold_WRDATA2_WRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
tsetup_WRDATA1_WRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
thold_WRDATA1_WRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
tsetup_WRDATA0_WRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
thold_WRDATA0_WRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
tsetup_WRAD4_WRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
thold_WRAD4_WRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
tsetup_WRAD3_WRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
thold_WRAD3_WRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
tsetup_WRAD2_WRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
thold_WRAD2_WRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
tsetup_WRAD1_WRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
thold_WRAD1_WRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
tsetup_WRAD0_WRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
thold_WRAD0_WRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
tpw_WRCLK_posedge        :VitalDelayType := 1.0 ns;
tpw_ADRCLK_posedge        :VitalDelayType := 1.0 ns;
tsetup_WEN_ADRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
thold_WEN_ADRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
tsetup_WRAD4_ADRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
thold_WRAD4_ADRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
tsetup_WRAD3_ADRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
thold_WRAD3_ADRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
tsetup_WRAD2_ADRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
thold_WRAD2_ADRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
tsetup_WRAD1_ADRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
thold_WRAD1_ADRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
tsetup_WRAD0_ADRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
thold_WRAD0_ADRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;
 
 
	TimingChecksOn : BOOLEAN := TRUE; 
	InstancePath : STRING := "*" 
            ); 
  PORT	( 
	WEN		: IN	std_logic ; 
	WRCLK		: IN	std_logic ; 
	ADRCLK		: IN	std_logic ; 
	OE		: IN	std_logic ; 
        WRDATA3         : INOUT std_logic := 'Z';
        WRDATA2         : INOUT std_logic := 'Z';
        WRDATA1         : INOUT std_logic := 'Z';
        WRDATA0         : INOUT std_logic := 'Z';
        WRAD4           : IN    std_logic;
        WRAD3           : IN    std_logic;
        WRAD2           : IN    std_logic;
        WRAD1           : IN    std_logic;
        WRAD0           : IN    std_logic
	); 
 
 
   ATTRIBUTE VITAL_LEVEL0 OF RB_MAR : ENTITY IS TRUE; 
 
END RB_MAR; 
 
----------------------------------------------------------------------- 
-- ARCHITECTURE declaration 
----------------------------------------------------------------------- 
ARCHITECTURE VITAL_VF OF RB_MAR IS 
 
    ATTRIBUTE VITAL_LEVEL1 OF VITAL_VF : ARCHITECTURE IS FALSE; 
 
	SIGNAL WEN_ipd		: std_logic := 'X'; 
	SIGNAL WRCLK_ipd		: std_logic := '0'; 
	SIGNAL ADRCLK_ipd		: std_logic := '0'; 
	SIGNAL WR_CLK		: std_logic := '0'; 
	SIGNAL ADR_CLK		: std_logic := '0'; 
	SIGNAL OE_ipd	: std_logic := 'X'; 
	SIGNAL DIN		: std_logic_vector(3 DOWNTO 0); 
	SIGNAL RD_ADD_W		: std_logic_vector(4 DOWNTO 0); 
	SIGNAL r_add_w		: std_logic_vector(4 DOWNTO 0); 
	SIGNAL WR_ADD		: std_logic_vector(4 DOWNTO 0); 
        SIGNAL WRDATA3_ipd      : std_logic := 'Z';
        SIGNAL WRDATA2_ipd      : std_logic := 'Z';
        SIGNAL WRDATA1_ipd      : std_logic := 'Z';
        SIGNAL WRDATA0_ipd      : std_logic := 'Z';
        SIGNAL WRAD4_ipd                : std_logic := '0';
        SIGNAL WRAD3_ipd                : std_logic := '0';
        SIGNAL WRAD2_ipd                : std_logic := '0';
        SIGNAL WRAD1_ipd                : std_logic := '0';
        SIGNAL WRAD0_ipd                : std_logic := '0';
	SIGNAL write_add	: std_logic_vector(4 DOWNTO 0); 
	SIGNAL data_out_w		: std_logic_vector(3 DOWNTO 0) := x_data; 
	SIGNAL output_delay	: time		:= 0 ns; 
	SIGNAL memory_array	: memory_array_typ; 
 
BEGIN 
    
  --------------------------------------------------------------------- 
  -- INPUT PATH DELAYs 
  --------------------------------------------------------------------- 
  WIREDELAY : BLOCK 
  BEGIN 
	VitalWireDelay (WEN_ipd,		WEN,		tipd_WEN); 
	VitalWireDelay (WRCLK_ipd,		WRCLK,		tipd_WRCLK); 
	VitalWireDelay (ADRCLK_ipd,		ADRCLK,		tipd_ADRCLK); 
	VitalWireDelay (OE_ipd,		OE,		tipd_OE); 
        VitalWireDelay (WRDATA0_ipd,    WRDATA0,        tipd_WRDATA0);
        VitalWireDelay (WRDATA1_ipd,    WRDATA1,        tipd_WRDATA1);
        VitalWireDelay (WRDATA2_ipd,    WRDATA2,        tipd_WRDATA2);
        VitalWireDelay (WRDATA3_ipd,    WRDATA3,        tipd_WRDATA3);
        VitalWireDelay (WRAD0_ipd,              WRAD0,          tipd_WRAD0);
        VitalWireDelay (WRAD1_ipd,              WRAD1,          tipd_WRAD1);
        VitalWireDelay (WRAD2_ipd,              WRAD2,          tipd_WRAD2);
        VitalWireDelay (WRAD3_ipd,              WRAD3,          tipd_WRAD3);
        VitalWireDelay (WRAD4_ipd,              WRAD4,          tipd_WRAD4); 
  END BLOCK; 
 
  --------------------------------------------------------------------- 
  -- Behavior Section 
  --------------------------------------------------------------------- 
 
  --------------------------------------------------------------------- 
  -- Wrapper Section 
  --------------------------------------------------------------------- 
 
   wrapper_latch_add_w : process(ADR_CLK)
   
   begin
      if (ADR_CLK = '1') then
           r_add_w(4) <= WRAD4_ipd;
           r_add_w(3) <= WRAD3_ipd;
           r_add_w(2) <= WRAD2_ipd;
           r_add_w(1) <= WRAD1_ipd;
           r_add_w(0) <= WRAD0_ipd;
      end if;

   end process;

   wrapper_read_add : process(r_add_w) 
 
   begin 
	RD_ADD_W <= r_add_w; 
   end process; 
 
   wrapper_write_add : process(WEN_ipd, WRAD4_ipd, WRAD3_ipd, WRAD2_ipd, WRAD1_ipd, WRAD0_ipd) 
 
   begin 
    if (WEN_ipd = '1') then 
        WR_ADD(4) <= WRAD4_ipd;
        WR_ADD(3) <= WRAD3_ipd;
        WR_ADD(2) <= WRAD2_ipd;
        WR_ADD(1) <= WRAD1_ipd;
        WR_ADD(0) <= WRAD0_ipd;
    else 
	WR_ADD <= x_add; 
    end if; 
 
   end process; 
 
   wrapper_write_clk : process(WEN_ipd, WRCLK_ipd) 
 
   begin 
    if (WEN_ipd = '1') then 
	WR_CLK <= WRCLK_ipd; 
    else 
	WR_CLK <= '0'; 
    end if; 
 
   end process; 

   wrapper_addr_clk : process(ADRCLK_ipd,WEN_ipd) 
 
   begin 
      if (WEN_ipd = '0') then
	ADR_CLK <= ADRCLK_ipd; 
      else
        ADR_CLK <= '0';
      end if;
    end process; 
 
   process(WR_CLK) 
 
    begin 
      if WR_CLK = '1' then 
        write_add(4) <= WRAD4_ipd;
        write_add(3) <= WRAD3_ipd;
        write_add(2) <= WRAD2_ipd;
        write_add(1) <= WRAD1_ipd;
        write_add(0) <= WRAD0_ipd;
      end if; 
 
   end process; 
 
   wrapper_write_data : process(WEN_ipd, WRDATA3_ipd, WRDATA2_ipd, WRDATA1_ipd, WRDATA0_ipd) 
 
   begin 
    if (WEN_ipd = '1') then 
        DIN(3) <= WRDATA3_ipd;
        DIN(2) <= WRDATA2_ipd;
        DIN(1) <= WRDATA1_ipd;
        DIN(0) <= WRDATA0_ipd;
    else 
	DIN <= x_data; 
    end if; 
 
   end process; 
 
 
  VITALBehavior : PROCESS ( WEN_ipd, WR_CLK, ADRCLK, ADR_CLK,  DIN, RD_ADD_W, WR_ADD ) 
 
 
   -- Temporary variables 
   VARIABLE tempaddr 		: integer := 0; 
   VARIABLE rd_address 	: integer := 0; 
   VARIABLE rd_viol_flag 	: X01 := '0'; 
 
   -- Timing Check results 
   VARIABLE Pviol_WRCLK			: std_logic := '0'; 
   VARIABLE PeriodData_WRCLK		: VitalPeriodDataType := VitalPeriodDataInit; 
   VARIABLE Pviol_ADRCLK			: std_logic := '0'; 
   VARIABLE PeriodData_ADRCLK		: VitalPeriodDataType := VitalPeriodDataInit; 
   VARIABLE Tviol_WR_ADD_stp_hld_0	: std_logic := '0'; 
   VARIABLE TimingData_WR_ADD_stp_hld_0	: VitalTimingDataType := VitalTimingDataInit; 
   VARIABLE Tviol_WR_ADD_stp_hld_1	: std_logic := '0'; 
   VARIABLE TimingData_WR_ADD_stp_hld_1	: VitalTimingDataType := VitalTimingDataInit; 
   VARIABLE Tviol_WR_ADD_stp_hld_2	: std_logic := '0'; 
   VARIABLE TimingData_WR_ADD_stp_hld_2	: VitalTimingDataType := VitalTimingDataInit; 
   VARIABLE Tviol_WR_ADD_stp_hld_3	: std_logic := '0'; 
   VARIABLE TimingData_WR_ADD_stp_hld_3	: VitalTimingDataType := VitalTimingDataInit; 
   VARIABLE Tviol_WR_ADD_stp_hld_4	: std_logic := '0'; 
   VARIABLE TimingData_WR_ADD_stp_hld_4	: VitalTimingDataType := VitalTimingDataInit; 
   VARIABLE Tviol_WR_DATA_stp_0		: std_logic := '0'; 
   VARIABLE TimingData_WR_DATA_stp_0	: VitalTimingDataType := VitalTimingDataInit; 
   VARIABLE Tviol_WR_DATA_stp_1		: std_logic := '0'; 
   VARIABLE TimingData_WR_DATA_stp_1	: VitalTimingDataType := VitalTimingDataInit; 
   VARIABLE Tviol_WR_DATA_stp_2		: std_logic := '0'; 
   VARIABLE TimingData_WR_DATA_stp_2	: VitalTimingDataType := VitalTimingDataInit; 
   VARIABLE Tviol_WR_DATA_stp_3		: std_logic := '0'; 
   VARIABLE TimingData_WR_DATA_stp_3	: VitalTimingDataType := VitalTimingDataInit; 
   VARIABLE Tviol_WR_DATA_hld_0		: std_logic := '0'; 
   VARIABLE TimingData_WR_DATA_hld_0	: VitalTimingDataType := VitalTimingDataInit; 
   VARIABLE Tviol_WR_DATA_hld_1		: std_logic := '0'; 
   VARIABLE TimingData_WR_DATA_hld_1	: VitalTimingDataType := VitalTimingDataInit; 
   VARIABLE Tviol_WR_DATA_hld_2		: std_logic := '0'; 
   VARIABLE TimingData_WR_DATA_hld_2	: VitalTimingDataType := VitalTimingDataInit; 
   VARIABLE Tviol_WR_DATA_hld_3		: std_logic := '0'; 
   VARIABLE TimingData_WR_DATA_hld_3	: VitalTimingDataType := VitalTimingDataInit; 
   VARIABLE Tviol_RD_ADD_stp_hld_0		: std_logic := '0'; 
   VARIABLE TimingData_RD_ADD_stp_hld_0	: VitalTimingDataType := VitalTimingDataInit; 
   VARIABLE Tviol_RD_ADD_stp_hld_1		: std_logic := '0'; 
   VARIABLE TimingData_RD_ADD_stp_hld_1	: VitalTimingDataType := VitalTimingDataInit; 
   VARIABLE Tviol_RD_ADD_stp_hld_2		: std_logic := '0'; 
   VARIABLE TimingData_RD_ADD_stp_hld_2	: VitalTimingDataType := VitalTimingDataInit; 
   VARIABLE Tviol_RD_ADD_stp_hld_3		: std_logic := '0'; 
   VARIABLE TimingData_RD_ADD_stp_hld_3	: VitalTimingDataType := VitalTimingDataInit; 
   VARIABLE Tviol_RD_ADD_stp_hld_4		: std_logic := '0'; 
   VARIABLE TimingData_RD_ADD_stp_hld_4	: VitalTimingDataType := VitalTimingDataInit; 
   VARIABLE Tviol_WEN_hld		: std_logic := '0'; 
   VARIABLE TimingData_WEN_hld		: VitalTimingDataType := VitalTimingDataInit; 
 
 
 
 BEGIN 
    ------------------------------------------------------------------- 
    -- Timing Check Section 
    ------------------------------------------------------------------- 
    IF (TimingChecksOn) THEN 
 
	VitalPeriodPulseCheck  (Pviol_WRCLK, 
				PeriodData_WRCLK, 
				WR_CLK, "WRCLK", 
				0.0 ns, 
				0.0 ns, 
				tpw_WRCLK_posedge, 
				0.0 ns, 
				True,
				InstancePath & "/RB_MAR", 
				TRUE, 
				TRUE, 
				WARNING ); 

	VitalPeriodPulseCheck  (Pviol_ADRCLK, 
				PeriodData_ADRCLK, 
				ADR_CLK, "ADRCLK", 
				0.0 ns, 
				0.0 ns, 
				tpw_ADRCLK_posedge, 
				0.0 ns, 
				True,
				InstancePath & "/RB_MAR", 
				TRUE, 
				TRUE, 
				WARNING ); 
 
        VitalSetupHoldCheck    (Tviol_WR_ADD_stp_hld_0,
                                TimingData_WR_ADD_stp_hld_0,
                                WR_ADD(0), "WRAD0",
                                0.0 ns,
                                WR_CLK, "WRCLK",
                                0.0 ns,
                                tsetup_WRAD0_WRCLK_noedge_posedge, tsetup_WRAD0_WRCLK_noedge_posedge,
                                thold_WRAD0_WRCLK_noedge_posedge, thold_WRAD0_WRCLK_noedge_posedge,
                                WEN_ipd = '1',
                                '/',
                                InstancePath & "/RB_MAR",
                                TRUE,
                                TRUE,
                                WARNING );

        VitalSetupHoldCheck    (Tviol_WR_ADD_stp_hld_1,
                                TimingData_WR_ADD_stp_hld_1,
                                WR_ADD(1), "WRAD1",
                                0.0 ns,
                                WR_CLK, "WRCLK",
                                0.0 ns,
                                tsetup_WRAD1_WRCLK_noedge_posedge, tsetup_WRAD1_WRCLK_noedge_posedge,
                                thold_WRAD1_WRCLK_noedge_posedge, thold_WRAD1_WRCLK_noedge_posedge,
                                WEN_ipd = '1',
                                '/',
                                InstancePath & "/RB_MAR",
                                TRUE,
                                TRUE,
                                WARNING );

        VitalSetupHoldCheck    (Tviol_WR_ADD_stp_hld_2,
                                TimingData_WR_ADD_stp_hld_2,
                                WR_ADD(2), "WRAD2",
                                0.0 ns,
                                WR_CLK, "WRCLK",
                                0.0 ns,
                                tsetup_WRAD2_WRCLK_noedge_posedge, tsetup_WRAD2_WRCLK_noedge_posedge,
                                thold_WRAD2_WRCLK_noedge_posedge, thold_WRAD2_WRCLK_noedge_posedge,
                                WEN_ipd = '1',
                                '/',
                                InstancePath & "/RB_MAR",
                                TRUE,
                                TRUE,
                                WARNING );
       VitalSetupHoldCheck    (Tviol_WR_ADD_stp_hld_3,
                                TimingData_WR_ADD_stp_hld_3,
                                WR_ADD(3), "WRAD3",
                                0.0 ns,
                                WR_CLK, "WRCLK",
                                0.0 ns,
                                tsetup_WRAD3_WRCLK_noedge_posedge, tsetup_WRAD3_WRCLK_noedge_posedge,
                                thold_WRAD3_WRCLK_noedge_posedge, thold_WRAD3_WRCLK_noedge_posedge,
                                WEN_ipd = '1',
                                '/',
                                InstancePath & "/RB_MAR",
                                TRUE,
                                TRUE,
                                WARNING );
  VitalSetupHoldCheck    (Tviol_WR_ADD_stp_hld_4,
                                TimingData_WR_ADD_stp_hld_4,
                                WR_ADD(4), "WRAD4",
                                0.0 ns,
                                WR_CLK, "WRCLK",
                                0.0 ns,
                                tsetup_WRAD4_WRCLK_noedge_posedge, tsetup_WRAD4_WRCLK_noedge_posedge,
                                thold_WRAD4_WRCLK_noedge_posedge, thold_WRAD4_WRCLK_noedge_posedge,
                                WEN_ipd = '1',
                                '/',
                                InstancePath & "/RB_MAR",
                                TRUE,
                                TRUE,
                                WARNING );

        VitalSetupHoldCheck    (Tviol_WR_DATA_stp_0,
                                TimingData_WR_DATA_stp_0,
                                DIN(0), "WRDATA0",
                                0.0 ns,
                                WR_CLK, "WRCLK",
                                0.0 ns,
                                tsetup_WRDATA0_WRCLK_noedge_posedge, tsetup_WRDATA0_WRCLK_noedge_posedge,
                                0.0 ns, 0.0 ns,
                                WEN_ipd = '1',
                                '/',
                                InstancePath & "/RB_MAR",
                                TRUE,
                                TRUE,
                                WARNING );

        VitalSetupHoldCheck    (Tviol_WR_DATA_stp_1,
                                TimingData_WR_DATA_stp_1,
                                DIN(1), "WRDATA1",
                                0.0 ns,
                                WR_CLK, "WRCLK",
                                0.0 ns,
                                tsetup_WRDATA1_WRCLK_noedge_posedge, tsetup_WRDATA1_WRCLK_noedge_posedge,
                                0.0 ns, 0.0 ns,
                                WEN_ipd = '1',
                                '/',
                                InstancePath & "/RB_MAR",
                                TRUE,
                                TRUE,
                                WARNING );

        VitalSetupHoldCheck    (Tviol_WR_DATA_stp_2,
                                TimingData_WR_DATA_stp_2,
                                DIN(2), "WRDATA2",
                                0.0 ns,
                                WR_CLK, "WRCLK",
                                0.0 ns,
                                tsetup_WRDATA2_WRCLK_noedge_posedge, tsetup_WRDATA2_WRCLK_noedge_posedge,
                                0.0 ns, 0.0 ns,
                                WEN_ipd = '1',
                                '/',
                                InstancePath & "/RB_MAR",
                                TRUE,
                                TRUE,
                                WARNING );
        VitalSetupHoldCheck    (Tviol_WR_DATA_stp_3,
                                TimingData_WR_DATA_stp_3,
                                DIN(3), "WRDATA3",
                                0.0 ns,
                                WR_CLK, "WRCLK",
                                0.0 ns,
                                tsetup_WRDATA3_WRCLK_noedge_posedge, tsetup_WRDATA3_WRCLK_noedge_posedge,
                                0.0 ns, 0.0 ns,
                                WEN_ipd = '1',
                                '/',
                                InstancePath & "/RB_MAR",
                                TRUE,
                                TRUE,
                                WARNING );

        VitalSetupHoldCheck    (Tviol_WR_DATA_hld_0,
                                TimingData_WR_DATA_hld_0,
                                DIN(0), "WRDATA0",
                                0.0 ns,
                                WR_CLK, "WRCLK",
                                0.0 ns,
                                0.0 ns, 0.0 ns,
                                thold_WRDATA0_WRCLK_noedge_posedge, thold_WRDATA0_WRCLK_noedge_posedge,
                                WEN_ipd = '1',
                                '/',
                                InstancePath & "/RB_MAR",
                                TRUE,
                                TRUE,
                                WARNING );

        VitalSetupHoldCheck    (Tviol_WR_DATA_hld_1,
                                TimingData_WR_DATA_hld_1,
                                DIN(1), "WRDATA1",
                                0.0 ns,
                                WR_CLK, "WRCLK",
                                0.0 ns,
                                0.0 ns, 0.0 ns,
                                thold_WRDATA1_WRCLK_noedge_posedge, thold_WRDATA1_WRCLK_noedge_posedge,
                                WEN_ipd = '1',
                                '/',
                                InstancePath & "/RB_MAR",
                                TRUE,
                                TRUE,
                                WARNING );

        VitalSetupHoldCheck    (Tviol_WR_DATA_hld_2,
                                TimingData_WR_DATA_hld_2,
                                DIN(2), "WRDATA2",
                                0.0 ns,
                                WR_CLK, "WRCLK",
                                0.0 ns,
                                0.0 ns, 0.0 ns,
                                thold_WRDATA2_WRCLK_noedge_posedge, thold_WRDATA2_WRCLK_noedge_posedge,
                                WEN_ipd = '1',
                                '/',
                                InstancePath & "/RB_MAR",
                                TRUE,
                                TRUE,
                                WARNING );
        VitalSetupHoldCheck    (Tviol_WR_DATA_hld_3,
                                TimingData_WR_DATA_hld_3,
                                DIN(3), "WRDATA3",
                                0.0 ns,
                                WR_CLK, "WRCLK",
                                0.0 ns,
                                0.0 ns, 0.0 ns,
                                thold_WRDATA3_WRCLK_noedge_posedge, thold_WRDATA3_WRCLK_noedge_posedge,
                                WEN_ipd = '1',
                                '/',
                                InstancePath & "/RB_MAR",
                                TRUE,
                                TRUE,
                                WARNING );
        VitalSetupHoldCheck    (Tviol_RD_ADD_stp_hld_0,
                                TimingData_RD_ADD_stp_hld_0,
                                WRAD0_ipd, "WRAD0",
                                0.0 ns,
                                ADRCLK_ipd, "ADRCLK",
                                0.0 ns,
                                tsetup_WRAD0_ADRCLK_noedge_posedge, tsetup_WRAD0_ADRCLK_noedge_posedge,
                                thold_WRAD0_ADRCLK_noedge_posedge, thold_WRAD0_ADRCLK_noedge_posedge,
                                True,
                                '/',
                                InstancePath & "/RB_MAR",
                                TRUE,
                                TRUE,
                                WARNING );

        VitalSetupHoldCheck    (Tviol_RD_ADD_stp_hld_1,
                                TimingData_RD_ADD_stp_hld_1,
                                WRAD1_ipd, "WRAD1",
                                0.0 ns,
                                ADRCLK_ipd, "ADRCLK",
                                0.0 ns,
                                tsetup_WRAD1_ADRCLK_noedge_posedge, tsetup_WRAD1_ADRCLK_noedge_posedge,
                                thold_WRAD1_ADRCLK_noedge_posedge, thold_WRAD1_ADRCLK_noedge_posedge,
                                True,
                                '/',
                                InstancePath & "/RB_MAR",
                                TRUE,
                                TRUE,
                                WARNING );

        VitalSetupHoldCheck    (Tviol_RD_ADD_stp_hld_2,
                                TimingData_RD_ADD_stp_hld_2,
                                WRAD2_ipd, "WRAD2",
                                0.0 ns,
                                ADRCLK_ipd, "ADRCLK",
                                0.0 ns,
                                tsetup_WRAD2_ADRCLK_noedge_posedge, tsetup_WRAD2_ADRCLK_noedge_posedge,
                                thold_WRAD2_ADRCLK_noedge_posedge, thold_WRAD2_ADRCLK_noedge_posedge,
                                True,
                                '/',
                                InstancePath & "/RB_MAR",
                                TRUE,
                                TRUE,
                                WARNING );

        VitalSetupHoldCheck    (Tviol_RD_ADD_stp_hld_3,
                                TimingData_RD_ADD_stp_hld_3,
                                WRAD3_ipd, "WRAD3",
                                0.0 ns,
                                ADRCLK_ipd, "ADRCLK",
                                0.0 ns,
                                tsetup_WRAD3_ADRCLK_noedge_posedge, tsetup_WRAD3_ADRCLK_noedge_posedge,
                                thold_WRAD3_ADRCLK_noedge_posedge, thold_WRAD3_ADRCLK_noedge_posedge,
                                True,
                                '/',
                                InstancePath & "/RB_MAR",
                                TRUE,
                                TRUE,
                                WARNING );
        VitalSetupHoldCheck    (Tviol_RD_ADD_stp_hld_4,
                                TimingData_RD_ADD_stp_hld_4,
                                WRAD4_ipd, "WRAD4",
                                0.0 ns,
                                ADRCLK_ipd, "ADRCLK",
                                0.0 ns,
                                tsetup_WRAD4_ADRCLK_noedge_posedge, tsetup_WRAD4_ADRCLK_noedge_posedge,
                                thold_WRAD4_ADRCLK_noedge_posedge, thold_WRAD4_ADRCLK_noedge_posedge,
                                True,
                                '/',
                                InstancePath & "/RB_MAR",
                                TRUE,
                                TRUE,
                                WARNING );

	VitalSetupHoldCheck    (Tviol_WEN_hld, 
				TimingData_WEN_hld, 
				WEN_ipd, "WEN", 
				0.0 ns, 
				ADR_CLK, "ADRCLK", 
				0.0 ns, 
				tsetup_WEN_ADRCLK_noedge_posedge, tsetup_WEN_ADRCLK_noedge_posedge,
				thold_WEN_ADRCLK_noedge_posedge, thold_WEN_ADRCLK_noedge_posedge,
				True, 
				'/', 
				InstancePath & "/RB_MAR", 
				TRUE, 
				TRUE, 
				WARNING ); 
 
    END IF; -- Timing Check Section 

 
 rd_viol_flag :=  (Tviol_RD_ADD_stp_hld_0 or Tviol_RD_ADD_stp_hld_1 or Tviol_RD_ADD_stp_hld_2 or Tviol_RD_ADD_stp_hld_3 or Tviol_RD_ADD_stp_hld_4 or Pviol_ADRCLK); 

 
 
 
    ------------------------------------------------------------------- 
    -- Functionality Section 
    ------------------------------------------------------------------- 
 
-- WRITE ADDRESS GOES XX 
 
    if ( WR_CLK'EVENT and WR_CLK = '1' and vecX(WR_ADD)) then 
 
        assert false 
        report "Illegal Address Input: Undefined  Address at the Read_Write Port." 
        severity note ; 
        memory_array <= (others => x_data); 
 
    end if; 
 
-- ADDRESS HOLD AND SETUP VIOLATION EFFECT 
 
    if( Tviol_WR_ADD_stp_hld_0 = 'X' or Tviol_WR_ADD_stp_hld_1 = 'X' or Tviol_WR_ADD_stp_hld_2 = 'X' or Tviol_WR_ADD_stp_hld_3 = 'X' or Tviol_WR_ADD_stp_hld_4 = 'X' ) then 
 
        memory_array <= (others => x_data); 
 
    else 
 
-- DATA SETUP AND HOLD VIOLATION EFFECT 
 
    if( Pviol_WRCLK = 'X' or Tviol_WR_DATA_hld_0 = 'X' or Tviol_WR_DATA_hld_1 = 'X' or Tviol_WR_DATA_hld_2 = 'X' or Tviol_WR_DATA_hld_3 = 'X' or Tviol_WEN_hld = 'X') then 
	tempaddr := vec2int(write_add); 
	memory_array(tempaddr) <= x_data; 
    end if; 
 
    if( Tviol_WR_DATA_stp_0 = 'X' or Tviol_WR_DATA_stp_1 = 'X' or Tviol_WR_DATA_stp_2 = 'X' or Tviol_WR_DATA_stp_3 = 'X') then 
	tempaddr := vec2int(WR_ADD); 
	memory_array(tempaddr) <= x_data; 
    end if; 
 
    end if; 
 
-- VALID MEMORY WRITE 
 
    if ( WR_CLK'EVENT and WR_CLK = '1' and not(vecX(WR_ADD)) and not(Tviol_WR_ADD_stp_hld_0 = 'X' or Tviol_WR_ADD_stp_hld_1 = 'X' or Tviol_WR_ADD_stp_hld_2 = 'X' or Tviol_WR_ADD_stp_hld_3 = 'X' or Tviol_WR_ADD_stp_hld_4 = 'X') and not( Pviol_WRCLK = 'X' or Tviol_WR_DATA_hld_0 = 'X' or Tviol_WR_DATA_hld_1 = 'X' or Tviol_WR_DATA_hld_2 = 'X' or Tviol_WR_DATA_hld_3 = 'X' or Tviol_WEN_hld = 'X') and not( Tviol_WR_DATA_stp_0 = 'X' or Tviol_WR_DATA_stp_1 = 'X' or Tviol_WR_DATA_stp_2 = 'X' or Tviol_WR_DATA_stp_3 = 'X')) then 
	tempaddr := vec2int(WR_ADD); 
	memory_array(tempaddr) <= DIN; 
    end if; 
 
    if WR_CLK'EVENT and WR_CLK /= WRCLK_ipd and WR_CLK'LAST_VALUE = '1' then 
	memory_array(tempaddr) <= x_data; 
    end if; 
 
 
-- READ CYCLE VIOLATION EFFECT 
 
-- VALID MEMORY READ 
 
   if( rd_viol_flag = 'X' or (OE_ipd'EVENT and OE_ipd = '1' and vecX(RD_ADD_W))) then
        data_out_w <= x_data;
    elsif
           
     (OE_ipd'EVENT and OE_ipd = '1' and not(rd_viol_flag = 'X') and not (vecX(RD_ADD_W))) then 
	rd_address := vec2int(RD_ADD_W); 
	data_out_w <= TRANSPORT memory_array(rd_address); 
    end if; 
 
 
-- VALID MEMORY READ 
 
  END PROCESS; 
 
    ------------------------------------------------------------------------------- 
    -- Temporary output signal should get assigned to the output signal. 
    ------------------------------------------------------------------------------- 
 
 
   PROCESS(data_out_w, WEN_ipd, OE_ipd, ADRCLK_ipd)

   VARIABLE GLITCH_DATA : VitalGlitchDataType;
   VARIABLE con : std_logic ;--:= '0';
    VARIABLE WEN_inv : std_logic ;--:= '0';
    VARIABLE WRDATA3_1 : std_logic := '0';--:= 'Z';
    VARIABLE WRDATA2_1 : std_logic := '0';--:= 'Z';
    VARIABLE WRDATA1_1 : std_logic := '0';--:= 'Z';
    VARIABLE WRDATA0_1 : std_logic := '0';--:= 'Z';

   BEGIN
       WEN_inv := VitalINV(WEN_ipd);
       con := VitalAND2(OE_ipd,WEN_inv);


      WRDATA3_1 := VITALBUFIF1(data_out_w(3),NOT(con));
      WRDATA2_1 := VITALBUFIF1(data_out_w(2),NOT(con));
      WRDATA1_1 := VITALBUFIF1(data_out_w(1),NOT(con));
      WRDATA0_1 := VITALBUFIF1(data_out_w(0),NOT(con));


      VitalPathDelay01Z ( WRDATA3, GLITCH_DATA, "WRDATA3", WRDATA3_1,
        Paths => (
        0 => ( ADRCLK_ipd'LAST_EVENT, VitalExtendToFillDelay(tpd_ADRCLK_WRDATA3), TRUE ),
        1 => ( OE_ipd'LAST_EVENT, VitalExtendToFillDelay(tpd_OE_WRDATA3), TRUE )),
        DefaultDelay=>VitalZeroDelay01Z,
        Mode=>VitalInertial,
        XON=>TRUE,
        MsgOn=>TRUE,
        MsgSeverity=>WARNING,
        OutputMap => "UX01ZWLH-");

      VitalPathDelay01Z ( WRDATA2, GLITCH_DATA, "WRDATA2", WRDATA2_1,
        Paths => (
        0 => ( ADRCLK_ipd'LAST_EVENT, VitalExtendToFillDelay(tpd_ADRCLK_WRDATA2), TRUE ),
        1 => ( OE_ipd'LAST_EVENT, VitalExtendToFillDelay(tpd_OE_WRDATA2), TRUE ) ),
        DefaultDelay=>VitalZeroDelay01Z,
        Mode=>VitalInertial,
        XON=>TRUE,
        MsgOn=>TRUE,
        MsgSeverity=>WARNING,
        OutputMap => "UX01ZWLH-");

      VitalPathDelay01Z ( WRDATA1, GLITCH_DATA, "WRDATA1", WRDATA1_1,
        Paths => (
        0 => ( ADRCLK_ipd'LAST_EVENT, VitalExtendToFillDelay(tpd_ADRCLK_WRDATA1), TRUE ),
        1 => ( OE_ipd'LAST_EVENT, VitalExtendToFillDelay(tpd_OE_WRDATA1), TRUE ) ),
        DefaultDelay=>VitalZeroDelay01Z,
        Mode=>VitalInertial,
        XON=>TRUE,
        MsgOn=>TRUE,
        MsgSeverity=>WARNING,
        OutputMap => "UX01ZWLH-");

       VitalPathDelay01Z ( WRDATA0, GLITCH_DATA, "WRDATA0", WRDATA0_1,
        Paths => (
        0 => ( ADRCLK_ipd'LAST_EVENT, VitalExtendToFillDelay(tpd_ADRCLK_WRDATA0), TRUE ),
        1 => ( OE_ipd'LAST_EVENT, VitalExtendToFillDelay(tpd_OE_WRDATA0), TRUE ) ),
        DefaultDelay=>VitalZeroDelay01Z,
        Mode=>VitalInertial,
        XON=>TRUE,
        MsgOn=>TRUE,
        MsgSeverity=>WARNING,
        OutputMap => "UX01ZWLH-");

END PROCESS;
 
 
END VITAL_VF; 
configuration CFG_RB_MAR_VITAL of RB_MAR is
        for VITAL_VF
        end for;
end CFG_RB_MAR_VITAL;
----------------------------------------------------------------------- 
 
-- VITAL model for RB_SAR 30.10 technology 
----------------------------------------------------------------------- 
 
LIBRARY IEEE; 
USE IEEE.std_logic_1164.ALL; 
USE IEEE.VITAL_timing.all; 
USE IEEE.VITAL_primitives.all; 
LIBRARY VF1; 
USE VF1.ALL; 
USE VF1.RAMPACK.ALL; 
 
----------------------------------------------------------------------- 
-- ENTITY declaration 
----------------------------------------------------------------------- 
 
ENTITY RB_SAR IS 
  GENERIC ( 
	tipd_WEN		: VitalDelayType01			:= (0.0 ns, 0.0 ns); 
	tipd_REN		: VitalDelayType01			:= (0.0 ns, 0.0 ns); 
	tipd_WCLK		: VitalDelayType01			:= (0.0 ns, 0.0 ns); 
	tipd_ADRCLK		: VitalDelayType01			:= (0.0 ns, 0.0 ns); 
        tipd_WDATA3             : VitalDelayType01                      := (0.0 ns, 0.0 ns);
        tipd_WDATA2             : VitalDelayType01                      := (0.0 ns, 0.0 ns);
        tipd_WDATA1             : VitalDelayType01                      := (0.0 ns, 0.0 ns);
        tipd_WDATA0             : VitalDelayType01                      := (0.0 ns, 0.0 ns);
        tipd_RAD4               : VitalDelayType01                      := (0.0 ns, 0.0 ns);
        tipd_RAD3               : VitalDelayType01                      := (0.0 ns, 0.0 ns);
        tipd_RAD2               : VitalDelayType01                      := (0.0 ns, 0.0 ns);
        tipd_RAD1               : VitalDelayType01                      := (0.0 ns, 0.0 ns);
        tipd_RAD0               : VitalDelayType01                      := (0.0 ns, 0.0 ns);
        tipd_WAD4               : VitalDelayType01                      := (0.0 ns, 0.0 ns);
        tipd_WAD3               : VitalDelayType01                      := (0.0 ns, 0.0 ns);
        tipd_WAD2               : VitalDelayType01                      := (0.0 ns, 0.0 ns);
        tipd_WAD1               : VitalDelayType01                      := (0.0 ns, 0.0 ns);
        tipd_WAD0               : VitalDelayType01                      := (0.0 ns, 0.0 ns);
 

 
tpd_ADRCLK_RDATA0         :VitalDelayType01 := (2.0 ns,2.0 ns);
tpd_ADRCLK_RDATA1         :VitalDelayType01 := (2.0 ns,2.0 ns);
tpd_ADRCLK_RDATA2         :VitalDelayType01 := (2.0 ns,2.0 ns);
tpd_ADRCLK_RDATA3         :VitalDelayType01 := (2.0 ns,2.0 ns);
tpd_REN_RDATA0         :VitalDelayType01 := (2.0 ns,2.0 ns);
tpd_REN_RDATA1         :VitalDelayType01 := (2.0 ns,2.0 ns);
tpd_REN_RDATA2         :VitalDelayType01 := (2.0 ns,2.0 ns);
tpd_REN_RDATA3         :VitalDelayType01 := (2.0 ns,2.0 ns);
tsetup_WDATA3_WCLK_noedge_posedge     :VitalDelayType := 1.0 ns;


thold_WDATA3_WCLK_noedge_posedge     :VitalDelayType := 1.0 ns;


tsetup_WDATA2_WCLK_noedge_posedge     :VitalDelayType := 1.0 ns;


thold_WDATA2_WCLK_noedge_posedge     :VitalDelayType := 1.0 ns;


tsetup_WDATA1_WCLK_noedge_posedge     :VitalDelayType := 1.0 ns;


thold_WDATA1_WCLK_noedge_posedge     :VitalDelayType := 1.0 ns;


tsetup_WDATA0_WCLK_noedge_posedge     :VitalDelayType := 1.0 ns;


thold_WDATA0_WCLK_noedge_posedge     :VitalDelayType := 1.0 ns;


tsetup_WAD4_WCLK_noedge_posedge     :VitalDelayType := 1.0 ns;


thold_WAD4_WCLK_noedge_posedge     :VitalDelayType := 1.0 ns;


tsetup_WAD3_WCLK_noedge_posedge     :VitalDelayType := 1.0 ns;


thold_WAD3_WCLK_noedge_posedge     :VitalDelayType := 1.0 ns;


tsetup_WAD2_WCLK_noedge_posedge     :VitalDelayType := 1.0 ns;


thold_WAD2_WCLK_noedge_posedge     :VitalDelayType := 1.0 ns;


tsetup_WAD1_WCLK_noedge_posedge     :VitalDelayType := 1.0 ns;


thold_WAD1_WCLK_noedge_posedge     :VitalDelayType := 1.0 ns;


tsetup_WAD0_WCLK_noedge_posedge     :VitalDelayType := 1.0 ns;


thold_WAD0_WCLK_noedge_posedge     :VitalDelayType := 1.0 ns;


tsetup_WEN_WCLK_noedge_posedge     :VitalDelayType := 1.0 ns;


thold_WEN_WCLK_noedge_posedge     :VitalDelayType := 1.0 ns;


tpw_WCLK_posedge        :VitalDelayType := 1.0 ns;

tpw_ADRCLK_posedge        :VitalDelayType := 1.0 ns;

tsetup_WEN_ADRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;


thold_WEN_ADRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;


tsetup_RAD4_ADRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;


thold_RAD4_ADRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;


tsetup_RAD3_ADRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;


thold_RAD3_ADRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;


tsetup_RAD2_ADRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;


thold_RAD2_ADRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;


tsetup_RAD1_ADRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;


thold_RAD1_ADRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;


tsetup_RAD0_ADRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;


thold_RAD0_ADRCLK_noedge_posedge     :VitalDelayType := 1.0 ns;




	TimingChecksOn : BOOLEAN := TRUE; 
	InstancePath : STRING := "*" 
            ); 
  PORT	( 
	WEN		: IN	std_logic ; 
	REN		: IN	std_logic ; 
	WCLK		: IN	std_logic ; 
	ADRCLK		: IN	std_logic ; 
        WDATA3          : IN    std_logic ;
        WDATA2          : IN    std_logic ;
        WDATA1          : IN    std_logic ;
        WDATA0          : IN    std_logic ;
        RDATA3          : OUT   std_logic ;
        RDATA2          : OUT   std_logic ;
        RDATA1          : OUT   std_logic ;
        RDATA0          : OUT   std_logic ;
        RAD4            : IN    std_logic ;
        RAD3            : IN    std_logic ;
        RAD2            : IN    std_logic ;
        RAD1            : IN    std_logic ;
        RAD0            : IN    std_logic ;
        WAD4            : IN    std_logic ;
        WAD3            : IN    std_logic ;
        WAD2            : IN    std_logic ;
        WAD1            : IN    std_logic ;
        WAD0            : IN    std_logic

	); 
 
 
   ATTRIBUTE VITAL_LEVEL0 OF RB_SAR : ENTITY IS TRUE; 
 
END RB_SAR; 
 
----------------------------------------------------------------------- 
-- ARCHITECTURE declaration 
----------------------------------------------------------------------- 
ARCHITECTURE VITAL_VF OF RB_SAR IS 
 
    ATTRIBUTE VITAL_LEVEL1 OF VITAL_VF : ARCHITECTURE IS FALSE; 
 
	SIGNAL WEN_ipd		: std_logic := 'X'; 
	SIGNAL REN_ipd		: std_logic := 'X'; 
	SIGNAL WCLK_ipd		: std_logic := '0'; 
	SIGNAL ADRCLK_ipd		: std_logic := '0'; 
	SIGNAL WR_CLK		: std_logic := '0'; 
        SIGNAL WDATA3_ipd       : std_logic := 'Z';
        SIGNAL WDATA2_ipd       : std_logic := 'Z';
        SIGNAL WDATA1_ipd       : std_logic := 'Z';
        SIGNAL WDATA0_ipd       : std_logic := 'Z';
        SIGNAL DIN              : std_logic_vector(3 DOWNTO 0);
        SIGNAL RAD4_ipd         : std_logic ;
        SIGNAL RAD3_ipd         : std_logic ;
        SIGNAL RAD2_ipd         : std_logic ;
        SIGNAL RAD1_ipd         : std_logic ;
        SIGNAL RAD0_ipd         : std_logic ;
        SIGNAL RD_ADD           : std_logic_vector(4 DOWNTO 0);
        SIGNAL WAD4_ipd         : std_logic ;
        SIGNAL WAD3_ipd         : std_logic ;
        SIGNAL WAD2_ipd         : std_logic ;
        SIGNAL WAD1_ipd         : std_logic ;
        SIGNAL WAD0_ipd         : std_logic ;
	SIGNAL r_add		: std_logic_vector(4 DOWNTO 0); 
	SIGNAL WR_ADD		: std_logic_vector(4 DOWNTO 0); 
	SIGNAL write_add	: std_logic_vector(4 DOWNTO 0); 
	SIGNAL data_out		: std_logic_vector(3 DOWNTO 0) := x_data; 
	SIGNAL output_delay	: time		:= 0 ns; 
	SIGNAL memory_array	: memory_array_typ; 
 
BEGIN 
    
  --------------------------------------------------------------------- 
  -- INPUT PATH DELAYs 
  --------------------------------------------------------------------- 
  WIREDELAY : BLOCK 
  BEGIN 
	VitalWireDelay (WEN_ipd,		WEN,		tipd_WEN); 
	VitalWireDelay (REN_ipd,		REN,		tipd_REN); 
	VitalWireDelay (WCLK_ipd,		WCLK,		tipd_WCLK); 
	VitalWireDelay (ADRCLK_ipd,		ADRCLK,		tipd_ADRCLK); 
        VitalWireDelay (WDATA0_ipd,             WDATA0,         tipd_WDATA0);
        VitalWireDelay (WDATA1_ipd,             WDATA1,         tipd_WDATA1);
        VitalWireDelay (WDATA2_ipd,             WDATA2,         tipd_WDATA2);
        VitalWireDelay (WDATA3_ipd,             WDATA3,         tipd_WDATA3);
        VitalWireDelay (RAD0_ipd,               RAD0,           tipd_RAD0);
        VitalWireDelay (RAD1_ipd,               RAD1,           tipd_RAD1);
        VitalWireDelay (RAD2_ipd,               RAD2,           tipd_RAD2);
        VitalWireDelay (RAD3_ipd,               RAD3,           tipd_RAD3);
        VitalWireDelay (RAD4_ipd,               RAD4,           tipd_RAD4);
        VitalWireDelay (WAD0_ipd,               WAD0,           tipd_WAD0);
        VitalWireDelay (WAD1_ipd,               WAD1,           tipd_WAD1);
        VitalWireDelay (WAD2_ipd,               WAD2,           tipd_WAD2);
        VitalWireDelay (WAD3_ipd,               WAD3,           tipd_WAD3);
        VitalWireDelay (WAD4_ipd,               WAD4,           tipd_WAD4);
 
  END BLOCK; 
 
  --------------------------------------------------------------------- 
  -- Behavior Section 
  --------------------------------------------------------------------- 
 
  --------------------------------------------------------------------- 
  -- Wrapper Section 
  --------------------------------------------------------------------- 
 
   wrapper_latch_add : process (ADRCLK_ipd)
   begin
     if (ADRCLK_ipd = '1') then
        r_add(4) <= RAD4_ipd;
        r_add(3) <= RAD3_ipd;
        r_add(2) <= RAD2_ipd;
        r_add(1) <= RAD1_ipd;
        r_add(0) <= RAD0_ipd;
     end if;
   end process;

   wrapper_read_add : process(r_add) 
 
   begin 
	RD_ADD <= r_add; 
 
   end process; 
 
 
  wrapper_write_add : process(WEN_ipd, WAD4_ipd, WAD3_ipd, WAD2_ipd, WAD1_ipd, WAD0_ipd)

   begin
    if (WEN_ipd = '1') then
        WR_ADD(4) <= WAD4_ipd;
        WR_ADD(3) <= WAD3_ipd;
        WR_ADD(2) <= WAD2_ipd;
        WR_ADD(1) <= WAD1_ipd;
        WR_ADD(0) <= WAD0_ipd;
    else
        WR_ADD <= x_add;
    end if;

   end process;

   wrapper_write_clk : process(WEN_ipd, WCLK_ipd) 
 
   begin 
    if (WEN_ipd = '1') then 
	WR_CLK <= WCLK_ipd; 
    else 
	WR_CLK <= '0'; 
    end if; 
 
   end process; 
 
    process(WR_CLK)

    begin
      if WR_CLK = '1' then
        write_add(4) <= WAD4_ipd;
        write_add(3) <= WAD3_ipd;
        write_add(2) <= WAD2_ipd;
        write_add(1) <= WAD1_ipd;
        write_add(0) <= WAD0_ipd;
      end if;

   end process;

   wrapper_write_data : process(WEN_ipd, WDATA3_ipd, WDATA2_ipd, WDATA1_ipd, WDATA0_ipd)

   begin
    if (WEN_ipd = '1') then
        DIN(3) <= WDATA3_ipd;
        DIN(2) <= WDATA2_ipd;
        DIN(1) <= WDATA1_ipd;
        DIN(0) <= WDATA0_ipd;
    else
        DIN <= x_data;
    end if;

   end process;
 
 
  VITALBehavior : PROCESS ( WEN_ipd, REN_ipd, WCLK_ipd, WR_CLK, RAD4_ipd, RAD3_ipd, RAD2_ipd, RAD1_ipd, RAD0_ipd, ADRCLK_ipd, DIN, RD_ADD, WR_ADD) 
 
 
   -- Temporary variables 
   VARIABLE tempaddr 		: integer := 0; 
   VARIABLE rd_address 		: integer := 0; 
   VARIABLE rd_viol_flag 	: X01 := '0'; 
 
   -- Timing Check results 
   VARIABLE Pviol_WCLK			: std_logic := '0'; 
   VARIABLE PeriodData_WCLK		: VitalPeriodDataType := VitalPeriodDataInit; 
   VARIABLE Pviol_ADRCLK			: std_logic := '0'; 
   VARIABLE PeriodData_ADRCLK		: VitalPeriodDataType := VitalPeriodDataInit; 
   VARIABLE Tviol_WR_ADD_stp_hld_0	: std_logic := '0'; 
   VARIABLE TimingData_WR_ADD_stp_hld_0	: VitalTimingDataType := VitalTimingDataInit; 
   VARIABLE Tviol_WR_ADD_stp_hld_1	: std_logic := '0'; 
   VARIABLE TimingData_WR_ADD_stp_hld_1	: VitalTimingDataType := VitalTimingDataInit; 
   VARIABLE Tviol_WR_ADD_stp_hld_2	: std_logic := '0'; 
   VARIABLE TimingData_WR_ADD_stp_hld_2	: VitalTimingDataType := VitalTimingDataInit; 
   VARIABLE Tviol_WR_ADD_stp_hld_3	: std_logic := '0'; 
   VARIABLE TimingData_WR_ADD_stp_hld_3	: VitalTimingDataType := VitalTimingDataInit; 
   VARIABLE Tviol_WR_ADD_stp_hld_4	: std_logic := '0'; 
   VARIABLE TimingData_WR_ADD_stp_hld_4	: VitalTimingDataType := VitalTimingDataInit; 
   VARIABLE Tviol_WR_DATA_stp_0		: std_logic := '0'; 
   VARIABLE TimingData_WR_DATA_stp_0	: VitalTimingDataType := VitalTimingDataInit; 
   VARIABLE Tviol_WR_DATA_stp_1		: std_logic := '0'; 
   VARIABLE TimingData_WR_DATA_stp_1	: VitalTimingDataType := VitalTimingDataInit; 
   VARIABLE Tviol_WR_DATA_stp_2		: std_logic := '0'; 
   VARIABLE TimingData_WR_DATA_stp_2	: VitalTimingDataType := VitalTimingDataInit; 
   VARIABLE Tviol_WR_DATA_stp_3		: std_logic := '0'; 
   VARIABLE TimingData_WR_DATA_stp_3	: VitalTimingDataType := VitalTimingDataInit; 
   VARIABLE Tviol_WEN_WCLK_stp_hld		: std_logic := '0'; 
   VARIABLE TimingData_WEN_WCLK_stp_hld		: VitalTimingDataType := VitalTimingDataInit; 
   VARIABLE Tviol_WEN_ADRCLK_stp_hld		: std_logic := '0'; 
   VARIABLE TimingData_WEN_ADRCLK_stp_hld		: VitalTimingDataType := VitalTimingDataInit; 
   VARIABLE Tviol_RD_ADD_stp_hld_0	: std_logic := '0'; 
   VARIABLE TimingData_RD_ADD_stp_hld_0	: VitalTimingDataType := VitalTimingDataInit; 
   VARIABLE Tviol_RD_ADD_stp_hld_1	: std_logic := '0'; 
   VARIABLE TimingData_RD_ADD_stp_hld_1	: VitalTimingDataType := VitalTimingDataInit; 
   VARIABLE Tviol_RD_ADD_stp_hld_2	: std_logic := '0'; 
   VARIABLE TimingData_RD_ADD_stp_hld_2	: VitalTimingDataType := VitalTimingDataInit; 
   VARIABLE Tviol_RD_ADD_stp_hld_3	: std_logic := '0'; 
   VARIABLE TimingData_RD_ADD_stp_hld_3	: VitalTimingDataType := VitalTimingDataInit; 
   VARIABLE Tviol_RD_ADD_stp_hld_4	: std_logic := '0'; 
   VARIABLE TimingData_RD_ADD_stp_hld_4	: VitalTimingDataType := VitalTimingDataInit; 
 
 
 
 BEGIN 
    ------------------------------------------------------------------- 
    -- Timing Check Section 
    ------------------------------------------------------------------- 
    IF (TimingChecksOn) THEN 
 
	VitalPeriodPulseCheck  (Pviol_WCLK, 
				PeriodData_WCLK, 
				WR_CLK, "WCLK", 
				0.0 ns, 
				0.0 ns, 
				tpw_WCLK_posedge, 
				0.0 ns, 
				TRUE,
				InstancePath & "/RB_SAR", 
				TRUE, 
				TRUE, 
				WARNING ); 

	VitalPeriodPulseCheck  (Pviol_ADRCLK, 
				PeriodData_ADRCLK, 
				ADRCLK, "ADRCLK", 
				0.0 ns, 
				0.0 ns, 
				tpw_ADRCLK_posedge, 
				0.0 ns, 
				True, 
				InstancePath & "/RB_SAR", 
				TRUE, 
				TRUE, 
				WARNING ); 
 
	VitalSetupHoldCheck    (Tviol_WR_ADD_stp_hld_0, 
				TimingData_WR_ADD_stp_hld_0, 
				WR_ADD(0), "WAD0", 
				0.0 ns, 
				WR_CLK, "WCLK", 
				0.0 ns, 
				tsetup_WAD0_WCLK_noedge_posedge, tsetup_WAD0_WCLK_noedge_posedge,  
				thold_WAD0_WCLK_noedge_posedge, thold_WAD0_WCLK_noedge_posedge, 
				WEN_ipd = '1', 
				'/', 
				InstancePath & "/RB_SAR", 
				TRUE, 
				TRUE, 
				WARNING ); 
 
	VitalSetupHoldCheck    (Tviol_WR_ADD_stp_hld_1, 
				TimingData_WR_ADD_stp_hld_1, 
				WR_ADD(1), "WAD1", 
				0.0 ns, 
				WR_CLK, "WCLK", 
				0.0 ns, 
				tsetup_WAD1_WCLK_noedge_posedge, tsetup_WAD1_WCLK_noedge_posedge,  
				thold_WAD1_WCLK_noedge_posedge, thold_WAD1_WCLK_noedge_posedge, 
				WEN_ipd = '1', 
				'/', 
				InstancePath & "/RB_SAR", 
				TRUE, 
				TRUE, 
				WARNING ); 
 
	VitalSetupHoldCheck    (Tviol_WR_ADD_stp_hld_2, 
				TimingData_WR_ADD_stp_hld_2, 
				WR_ADD(2), "WAD2", 
				0.0 ns, 
				WR_CLK, "WCLK", 
				0.0 ns, 
				tsetup_WAD2_WCLK_noedge_posedge, tsetup_WAD2_WCLK_noedge_posedge,  
				thold_WAD2_WCLK_noedge_posedge, thold_WAD2_WCLK_noedge_posedge, 
				WEN_ipd = '1', 
				'/', 
				InstancePath & "/RB_SAR", 
				TRUE, 
				TRUE, 
				WARNING ); 
 
	VitalSetupHoldCheck    (Tviol_WR_ADD_stp_hld_3, 
				TimingData_WR_ADD_stp_hld_3, 
				WR_ADD(3), "WAD3", 
				0.0 ns, 
				WR_CLK, "WCLK", 
				0.0 ns, 
				tsetup_WAD3_WCLK_noedge_posedge, tsetup_WAD3_WCLK_noedge_posedge,  
				thold_WAD3_WCLK_noedge_posedge, thold_WAD3_WCLK_noedge_posedge, 
				WEN_ipd = '1', 
				'/', 
				InstancePath & "/RB_SAR", 
				TRUE, 
				TRUE, 
				WARNING ); 
 
	VitalSetupHoldCheck    (Tviol_WR_ADD_stp_hld_4, 
				TimingData_WR_ADD_stp_hld_4, 
				WR_ADD(4), "WAD4", 
				0.0 ns, 
				WR_CLK, "WCLK", 
				0.0 ns, 
				tsetup_WAD4_WCLK_noedge_posedge, tsetup_WAD4_WCLK_noedge_posedge,  
				thold_WAD4_WCLK_noedge_posedge, thold_WAD4_WCLK_noedge_posedge, 
				WEN_ipd = '1', 
				'/', 
				InstancePath & "/RB_SAR", 
				TRUE, 
				TRUE, 
				WARNING ); 
 
	VitalSetupHoldCheck    (Tviol_WR_DATA_stp_0, 
				TimingData_WR_DATA_stp_0, 
				DIN(0), "WDATA0", 
				0.0 ns, 
				WR_CLK, "WCLK", 
				0.0 ns, 
				tsetup_WDATA0_WCLK_noedge_posedge, tsetup_WDATA0_WCLK_noedge_posedge,  
				thold_WDATA0_WCLK_noedge_posedge, thold_WDATA0_WCLK_noedge_posedge,  
				WEN_ipd = '1', 
				'/', 
				InstancePath & "/RB_SAR", 
				TRUE, 
				TRUE, 
				WARNING ); 
 
	VitalSetupHoldCheck    (Tviol_WR_DATA_stp_1, 
				TimingData_WR_DATA_stp_1, 
				DIN(1), "WDATA1", 
				0.0 ns, 
				WR_CLK, "WCLK", 
				0.0 ns, 
				tsetup_WDATA1_WCLK_noedge_posedge, tsetup_WDATA1_WCLK_noedge_posedge,  
				thold_WDATA1_WCLK_noedge_posedge, thold_WDATA1_WCLK_noedge_posedge,  
				WEN_ipd = '1', 
				'/', 
				InstancePath & "/RB_SAR", 
				TRUE, 
				TRUE, 
				WARNING ); 
 
	VitalSetupHoldCheck    (Tviol_WR_DATA_stp_2, 
				TimingData_WR_DATA_stp_2, 
				DIN(2), "WDATA2", 
				0.0 ns, 
				WR_CLK, "WCLK", 
				0.0 ns, 
				tsetup_WDATA2_WCLK_noedge_posedge, tsetup_WDATA2_WCLK_noedge_posedge,  
				thold_WDATA2_WCLK_noedge_posedge, thold_WDATA2_WCLK_noedge_posedge,  
				WEN_ipd = '1', 
				'/', 
				InstancePath & "/RB_SAR", 
				TRUE, 
				TRUE, 
				WARNING ); 
 
	VitalSetupHoldCheck    (Tviol_WR_DATA_stp_3, 
				TimingData_WR_DATA_stp_3, 
				DIN(3), "WDATA3", 
				0.0 ns, 
				WR_CLK, "WCLK", 
				0.0 ns, 
				tsetup_WDATA3_WCLK_noedge_posedge, tsetup_WDATA3_WCLK_noedge_posedge,  
				thold_WDATA3_WCLK_noedge_posedge, thold_WDATA3_WCLK_noedge_posedge,  
				WEN_ipd = '1', 
				'/', 
				InstancePath & "/RB_SAR", 
				TRUE, 
				TRUE, 
				WARNING ); 
 

        VitalSetupHoldCheck    (Tviol_RD_ADD_stp_hld_0,
                                TimingData_RD_ADD_stp_hld_0,
                                RAD0_ipd, "RAD0",
                                0.0 ns,
                                ADRCLK_ipd, "ADRCLK",
                                0.0 ns,
                                tsetup_RAD0_ADRCLK_noedge_posedge, tsetup_RAD0_ADRCLK_noedge_posedge,
                                thold_RAD0_ADRCLK_noedge_posedge, thold_RAD0_ADRCLK_noedge_posedge,
                                True,
                                '/',
                                InstancePath & "/RB_SAR",
                                TRUE,
                                TRUE,
                                WARNING );

        VitalSetupHoldCheck    (Tviol_RD_ADD_stp_hld_1,
                                TimingData_RD_ADD_stp_hld_1,
                                RAD1_ipd, "RAD1",
                                0.0 ns,
                                ADRCLK, "ADRCLK",
                                0.0 ns,
                                tsetup_RAD1_ADRCLK_noedge_posedge, tsetup_RAD1_ADRCLK_noedge_posedge,
                                thold_RAD1_ADRCLK_noedge_posedge, thold_RAD1_ADRCLK_noedge_posedge,
                                True,
                                '/',
                                InstancePath & "/RB_SAR",
                                TRUE,
                                TRUE,
                                WARNING );

        VitalSetupHoldCheck    (Tviol_RD_ADD_stp_hld_2,
                                TimingData_RD_ADD_stp_hld_2,
                                RAD2_ipd, "RAD2",
                                0.0 ns,
                                ADRCLK_ipd, "ADRCLK",
                                0.0 ns,
                                tsetup_RAD2_ADRCLK_noedge_posedge, tsetup_RAD2_ADRCLK_noedge_posedge,
                                thold_RAD2_ADRCLK_noedge_posedge, thold_RAD2_ADRCLK_noedge_posedge,
                                True,
                                '/',
                                InstancePath & "/RB_SAR",
                                TRUE,
                                TRUE,
                                WARNING );

        VitalSetupHoldCheck    (Tviol_RD_ADD_stp_hld_3,
                                TimingData_RD_ADD_stp_hld_3,
                                RAD3_ipd, "RAD3",
                                0.0 ns,
                                ADRCLK_ipd, "ADRCLK",
                                0.0 ns,
                                tsetup_RAD3_ADRCLK_noedge_posedge, tsetup_RAD3_ADRCLK_noedge_posedge,
                                thold_RAD3_ADRCLK_noedge_posedge, thold_RAD3_ADRCLK_noedge_posedge,
                                True,
                                '/',
                                InstancePath & "/RB_SAR",
                                TRUE,
                                TRUE,
                                WARNING );

        VitalSetupHoldCheck    (Tviol_RD_ADD_stp_hld_4,
                                TimingData_RD_ADD_stp_hld_4,
                                RAD4_ipd, "RAD4",
                                0.0 ns,
                                ADRCLK, "ADRCLK",
                                0.0 ns,
                                tsetup_RAD4_ADRCLK_noedge_posedge, tsetup_RAD4_ADRCLK_noedge_posedge,
                                thold_RAD4_ADRCLK_noedge_posedge, thold_RAD4_ADRCLK_noedge_posedge,
                                True,
                                '/',
                                InstancePath & "/RB_SAR",
                                TRUE,
                                TRUE,
                                WARNING );

        VitalSetupHoldCheck    (Tviol_WEN_WCLK_stp_hld,
                                TimingData_WEN_WCLK_stp_hld,
                                WEN, "WEN",
                                0.0 ns,
                                WCLK_ipd, "WCLK",
                                0.0 ns,
                                tsetup_WEN_WCLK_noedge_posedge, tsetup_WEN_WCLK_noedge_posedge,
                                thold_WEN_WCLK_noedge_posedge, thold_WEN_WCLK_noedge_posedge,
                                True,
                                '/',
                                InstancePath & "/RB_SAR",
                                TRUE,
                                TRUE,
                                WARNING );

        VitalSetupHoldCheck    (Tviol_WEN_ADRCLK_stp_hld,
                                TimingData_WEN_ADRCLK_stp_hld,
                                WEN, "WEN",
                                0.0 ns,
                                ADRCLK_ipd, "ADRCLK",
                                0.0 ns,
                                tsetup_WEN_ADRCLK_noedge_posedge, tsetup_WEN_ADRCLK_noedge_posedge,
                                thold_WEN_ADRCLK_noedge_posedge, thold_WEN_ADRCLK_noedge_posedge,
                                True,
                                '/',
                                InstancePath & "/RB_SAR",
                                TRUE,
                                TRUE,
                                WARNING );
 
    END IF; -- Timing Check Section 
 
 rd_viol_flag :=  (Tviol_RD_ADD_stp_hld_0 or Tviol_RD_ADD_stp_hld_1 or Tviol_RD_ADD_stp_hld_2 or Tviol_RD_ADD_stp_hld_3 or Tviol_RD_ADD_stp_hld_4 or Pviol_ADRCLK ); 
 
 
 
    ------------------------------------------------------------------- 
    -- Functionality Section 
    ------------------------------------------------------------------- 
 
-- WRITE ADDRESS GOES XX 
 
    if ( WR_CLK'EVENT and WR_CLK = '1' and vecX(WR_ADD)) then 
 
        assert false 
        report "Illegal Address Input: Undefined  Address at the Read_Write Port." 
        severity note ; 
        memory_array <= (others => x_data); 
 
    end if; 
 
-- ADDRESS HOLD AND SETUP VIOLATION EFFECT 
 
    if( Tviol_WR_ADD_stp_hld_0 = 'X' or Tviol_WR_ADD_stp_hld_1 = 'X' or Tviol_WR_ADD_stp_hld_2 = 'X' or Tviol_WR_ADD_stp_hld_3 = 'X' or Tviol_WR_ADD_stp_hld_4 = 'X' ) then 
 
        memory_array <= (others => x_data); 
 
    else 
 
-- DATA SETUP AND HOLD VIOLATION EFFECT 
 
 
    if( Pviol_WCLK = 'X' or Tviol_WR_DATA_stp_0 = 'X' or Tviol_WR_DATA_stp_1 = 'X' or Tviol_WR_DATA_stp_2 = 'X' or Tviol_WR_DATA_stp_3 = 'X') then 
	tempaddr := vec2int(WR_ADD); 
	memory_array(tempaddr) <= x_data; 
    end if; 
 
    end if; 
 
-- VALID MEMORY WRITE 
 
    if ( WR_CLK'EVENT and WR_CLK = '1' and not(vecX(WR_ADD)) and not(Tviol_WR_ADD_stp_hld_0 = 'X' or Tviol_WR_ADD_stp_hld_1 = 'X' or Tviol_WR_ADD_stp_hld_2 = 'X' or Tviol_WR_ADD_stp_hld_3 = 'X' or Tviol_WR_ADD_stp_hld_4 = 'X') and not(Tviol_WEN_WCLK_stp_hld = 'X') and not( Pviol_WCLK = 'X' or Tviol_WR_DATA_stp_0 = 'X' or Tviol_WR_DATA_stp_1 = 'X' or Tviol_WR_DATA_stp_2 = 'X' or Tviol_WR_DATA_stp_3 = 'X')) then 
	tempaddr := vec2int(WR_ADD); 
	memory_array(tempaddr) <= DIN; 
    end if; 
 
    if WR_CLK'EVENT and WR_CLK /= WCLK_ipd and WR_CLK'LAST_VALUE = '1' then 
	memory_array(tempaddr) <= x_data; 
    end if; 
 
 
-- READ CYCLE VIOLATION EFFECT 
 
    if( rd_viol_flag = 'X'  or (REN_ipd'EVENT  AND REN_ipd = '1'  and vecX(RD_ADD))) then 
	--output_delay <= 0 ns; 
	data_out <= x_data; 
    elsif 
 
-- VALID MEMORY READ 
 
 
     (((ADRCLK_ipd'EVENT and ADRCLK_ipd='1') or (REN_ipd'EVENT  and REN_ipd = '1'))  and not(rd_viol_flag = 'X') and not (vecX(RD_ADD))) then 
	rd_address := vec2int(RD_ADD); 
	--output_delay <= tpd_RAD_RDATA_X(0); 
	--data_out <= TRANSPORT x_data; 
	data_out <=  memory_array(rd_address); 
    end if; 
 
 
  END PROCESS; 
 
    ------------------------------------------------------------------------------- 
    -- Temporary output signal should get assigned to the output signal. 
    ------------------------------------------------------------------------------- 
 
 PROCESS(data_out, ADRCLK_ipd, REN_ipd)

   VARIABLE RDATA0_1 : std_logic := 'X';
   VARIABLE RDATA1_1 : std_logic := 'X';
   VARIABLE RDATA2_1 : std_logic := 'X';
   VARIABLE RDATA3_1 : std_logic := 'X';
   VARIABLE GLITCH_DATA : VitalGlitchDataType;
  BEGIN

    RDATA0_1 := VitalBUF(data_out(0));    --- Is this Vital level0 compliant
    RDATA1_1 := VitalBUF(data_out(1));
    RDATA2_1 := VitalBUF(data_out(2));
    RDATA3_1 := VitalBUF(data_out(3));

      VitalPathDelay01 ( RDATA3, GLITCH_DATA, "RDATA3", RDATA3_1,
        Paths => (
        0 => ( ADRCLK_ipd'LAST_EVENT, tpd_ADRCLK_RDATA3, TRUE ),
        1 => ( REN_ipd'LAST_EVENT, tpd_REN_RDATA3, TRUE ) ),
        DefaultDelay=>VitalZeroDelay01,
        Mode=>VitalInertial,
        XON=>TRUE,
        MsgOn=>TRUE,
        MsgSeverity=>WARNING );

      VitalPathDelay01 ( RDATA2, GLITCH_DATA, "RDATA2", RDATA2_1,
        Paths => (
        0 => ( ADRCLK_ipd'LAST_EVENT, tpd_ADRCLK_RDATA2, TRUE ),
        1 => ( REN_ipd'LAST_EVENT, tpd_REN_RDATA2, TRUE ) ),
        DefaultDelay=>VitalZeroDelay01,
        Mode=>VitalInertial,
        XON=>TRUE,
        MsgOn=>TRUE,
        MsgSeverity=>WARNING );

      VitalPathDelay01 ( RDATA1, GLITCH_DATA, "RDATA1", RDATA1_1,
        Paths => (
        0 => ( ADRCLK_ipd'LAST_EVENT, tpd_ADRCLK_RDATA1, TRUE ),
        1 => ( REN_ipd'LAST_EVENT, tpd_REN_RDATA1, TRUE ) ),
        DefaultDelay=>VitalZeroDelay01,
        Mode=>VitalInertial,
        XON=>TRUE,
        MsgOn=>TRUE,
        MsgSeverity=>WARNING );

      VitalPathDelay01 ( RDATA0, GLITCH_DATA, "RDATA0", RDATA0_1,
        Paths => (
        0 => ( ADRCLK_ipd'LAST_EVENT, tpd_ADRCLK_RDATA0, TRUE ),
        1 => ( REN_ipd'LAST_EVENT, tpd_REN_RDATA0, TRUE ) ),
        DefaultDelay=>VitalZeroDelay01,
        Mode=>VitalInertial,
        XON=>TRUE,
        MsgOn=>TRUE,
        MsgSeverity=>WARNING );

END PROCESS;

 
END VITAL_VF; 
configuration CFG_RB_SAR_VITAL of RB_SAR is
        for VITAL_VF
        end for;
end CFG_RB_SAR_VITAL;
----------------------------------------------------------------------- 
 
-----------------------------------------------------------------------
-- VITAL model for R_DA 30.10 technology
-----------------------------------------------------------------------

LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.VITAL_timing.all;
USE IEEE.std_logic_textio.all;
USE IEEE.VITAL_primitives.all;
LIBRARY std;
USE std.textio.all;
LIBRARY VF1;
USE VF1.ALL;
USE VF1.RAMPACK.ALL;

-----------------------------------------------------------------------
-- ENTITY declaration
-----------------------------------------------------------------------

ENTITY R_DA IS
  GENERIC (
	tipd_REN		: VitalDelayType01			:= (0.0 ns, 0.0 ns);
	tipd_OE		: VitalDelayType01			:= (0.0 ns, 0.0 ns);
	tipd_RAD14		: VitalDelayType01	:= (0.0 ns, 0.0 ns);
	tipd_RAD13		: VitalDelayType01	:= (0.0 ns, 0.0 ns);
	tipd_RAD12		: VitalDelayType01	:= (0.0 ns, 0.0 ns);
	tipd_RAD11		: VitalDelayType01	:= (0.0 ns, 0.0 ns);
	tipd_RAD10		: VitalDelayType01	:= (0.0 ns, 0.0 ns);
	tipd_RAD24		: VitalDelayType01	:= (0.0 ns, 0.0 ns);
	tipd_RAD23		: VitalDelayType01	:= (0.0 ns, 0.0 ns);
	tipd_RAD22		: VitalDelayType01	:= (0.0 ns, 0.0 ns);
	tipd_RAD21		: VitalDelayType01	:= (0.0 ns, 0.0 ns);
	tipd_RAD20		: VitalDelayType01	:= (0.0 ns, 0.0 ns);


	tpd_RAD14_RDATA13					: VitalDelayType01 := (2 ns,2 ns);
	tpd_RAD13_RDATA13					: VitalDelayType01 := (2 ns,2 ns);
	tpd_RAD12_RDATA13					: VitalDelayType01 := (2 ns,2 ns);
	tpd_RAD11_RDATA13					: VitalDelayType01 := (2 ns,2 ns);
	tpd_RAD10_RDATA13					: VitalDelayType01 := (2 ns,2 ns);
	tpd_RAD14_RDATA12					: VitalDelayType01 := (2 ns,2 ns);
	tpd_RAD13_RDATA12					: VitalDelayType01 := (2 ns,2 ns);
	tpd_RAD12_RDATA12					: VitalDelayType01 := (2 ns,2 ns);
	tpd_RAD11_RDATA12					: VitalDelayType01 := (2 ns,2 ns);
	tpd_RAD10_RDATA12					: VitalDelayType01 := (2 ns,2 ns);
	tpd_RAD14_RDATA11					: VitalDelayType01 := (2 ns,2 ns);
	tpd_RAD13_RDATA11					: VitalDelayType01 := (2 ns,2 ns);
	tpd_RAD12_RDATA11					: VitalDelayType01 := (2 ns,2 ns);
	tpd_RAD11_RDATA11					: VitalDelayType01 := (2 ns,2 ns);
	tpd_RAD10_RDATA11					: VitalDelayType01 := (2 ns,2 ns);
	tpd_RAD14_RDATA10					: VitalDelayType01 := (2 ns,2 ns);
	tpd_RAD13_RDATA10					: VitalDelayType01 := (2 ns,2 ns);
	tpd_RAD12_RDATA10					: VitalDelayType01 := (2 ns,2 ns);
	tpd_RAD11_RDATA10					: VitalDelayType01 := (2 ns,2 ns);
	tpd_RAD10_RDATA10					: VitalDelayType01 := (2 ns,2 ns);

	tpd_RAD24_RDATA23					: VitalDelayType01 := (2 ns,2 ns);
	tpd_RAD23_RDATA23					: VitalDelayType01 := (2 ns,2 ns);
	tpd_RAD22_RDATA23					: VitalDelayType01 := (2 ns,2 ns);
	tpd_RAD21_RDATA23					: VitalDelayType01 := (2 ns,2 ns);
	tpd_RAD20_RDATA23					: VitalDelayType01 := (2 ns,2 ns);
	tpd_RAD24_RDATA22					: VitalDelayType01 := (2 ns,2 ns);
	tpd_RAD23_RDATA22					: VitalDelayType01 := (2 ns,2 ns);
	tpd_RAD22_RDATA22					: VitalDelayType01 := (2 ns,2 ns);
	tpd_RAD21_RDATA22					: VitalDelayType01 := (2 ns,2 ns);
	tpd_RAD20_RDATA22					: VitalDelayType01 := (2 ns,2 ns);
	tpd_RAD24_RDATA21					: VitalDelayType01 := (2 ns,2 ns);
	tpd_RAD23_RDATA21					: VitalDelayType01 := (2 ns,2 ns);
	tpd_RAD22_RDATA21					: VitalDelayType01 := (2 ns,2 ns);
	tpd_RAD21_RDATA21					: VitalDelayType01 := (2 ns,2 ns);
	tpd_RAD20_RDATA21					: VitalDelayType01 := (2 ns,2 ns);
	tpd_RAD24_RDATA20					: VitalDelayType01 := (2 ns,2 ns);
	tpd_RAD23_RDATA20					: VitalDelayType01 := (2 ns,2 ns);
	tpd_RAD22_RDATA20					: VitalDelayType01 := (2 ns,2 ns);
	tpd_RAD21_RDATA20					: VitalDelayType01 := (2 ns,2 ns);
	tpd_RAD20_RDATA20					: VitalDelayType01 := (2 ns,2 ns);

	tpd_OE_RDATA23					: VitalDelayType01 := (2 ns,2 ns);
	tpd_OE_RDATA22					: VitalDelayType01 := (2 ns,2 ns);
	tpd_OE_RDATA21					: VitalDelayType01 := (2 ns,2 ns);
	tpd_OE_RDATA20					: VitalDelayType01 := (2 ns,2 ns);

	TimingChecksOn : BOOLEAN := TRUE;
	InstancePath : STRING := "*"
            );
  PORT	(
	REN		: IN	std_logic ;
	OE		: IN	std_logic ;
	RDATA23	        : OUT	std_logic := 'X';
	RDATA22	        : OUT	std_logic := 'X';
	RDATA21	        : OUT	std_logic := 'X';
	RDATA20	        : OUT	std_logic := 'X';
	RDATA13	        : OUT	std_logic := 'X';
	RDATA12	        : OUT	std_logic := 'X';
	RDATA11	        : OUT	std_logic := 'X';
	RDATA10	        : OUT	std_logic := 'X';
	RAD14		: IN	std_logic ;
	RAD13		: IN	std_logic ;
	RAD12		: IN	std_logic ;
	RAD11		: IN	std_logic ;
	RAD10		: IN	std_logic ;
	RAD24		: IN	std_logic ;
	RAD23		: IN	std_logic ;
	RAD22		: IN	std_logic ;
	RAD21		: IN	std_logic ;
	RAD20		: IN	std_logic 
	);


   ATTRIBUTE VITAL_LEVEL0 OF R_DA : ENTITY IS TRUE;

END R_DA;

-----------------------------------------------------------------------
-- ARCHITECTURE declaration
-----------------------------------------------------------------------
ARCHITECTURE VITAL_VF OF R_DA IS

    ATTRIBUTE VITAL_LEVEL1 OF VITAL_VF : ARCHITECTURE IS FALSE;

	file STF : text is in "rom_data";
	SIGNAL REN_ipd		: std_logic := 'X';
	SIGNAL OE_ipd	: std_logic := 'X';
	SIGNAL RAD14_ipd		: std_logic ;
	SIGNAL RAD13_ipd		: std_logic ;
	SIGNAL RAD12_ipd		: std_logic ;
	SIGNAL RAD11_ipd		: std_logic ;
	SIGNAL RAD10_ipd		: std_logic ;
	SIGNAL RD_ADD		: std_logic_vector(4 DOWNTO 0);
	SIGNAL RD_ADD2		: std_logic_vector(4 DOWNTO 0);
	SIGNAL RAD24_ipd		: std_logic ;
	SIGNAL RAD23_ipd		: std_logic ;
	SIGNAL RAD22_ipd		: std_logic ;
	SIGNAL RAD21_ipd		: std_logic ;
	SIGNAL RAD20_ipd		: std_logic ;
	SIGNAL data_out		: std_logic_vector(3 DOWNTO 0) := x_data;
	SIGNAL data_out_w	: std_logic_vector(3 DOWNTO 0) := x_data;
	SIGNAL output_delay	: time		:= 0 ns;
	SIGNAL output_delay_w	: time		:= 0 ns;
	SIGNAL memory_array	: memory_array_typ;

BEGIN
   
  ---------------------------------------------------------------------
  -- INPUT PATH DELAYs
  ---------------------------------------------------------------------
  WIREDELAY : BLOCK
  BEGIN
	VitalWireDelay (REN_ipd,		REN,		tipd_REN);
	VitalWireDelay (OE_ipd,		OE,		tipd_OE);
	VitalWireDelay (RAD10_ipd,		RAD10,		tipd_RAD10);
	VitalWireDelay (RAD11_ipd,		RAD11,		tipd_RAD11);
	VitalWireDelay (RAD12_ipd,		RAD12,		tipd_RAD12);
	VitalWireDelay (RAD13_ipd,		RAD13,		tipd_RAD13);
	VitalWireDelay (RAD14_ipd,		RAD14,		tipd_RAD14);
	VitalWireDelay (RAD20_ipd,		RAD20,	tipd_RAD20);
	VitalWireDelay (RAD21_ipd,		RAD21,	tipd_RAD21);
	VitalWireDelay (RAD22_ipd,		RAD22,	tipd_RAD22);
	VitalWireDelay (RAD23_ipd,		RAD23,	tipd_RAD23);
	VitalWireDelay (RAD24_ipd,		RAD24,	tipd_RAD24);

  END BLOCK;

  ---------------------------------------------------------------------
  -- Behavior Section
  ---------------------------------------------------------------------

  ---------------------------------------------------------------------
  -- Wrapper Section
  ---------------------------------------------------------------------

   wrapper_read_add : process(REN_ipd, RAD24_ipd, RAD23_ipd, RAD22_ipd, RAD21_ipd, RAD20_ipd, RAD14_ipd, RAD13_ipd, RAD12_ipd, RAD11_ipd, RAD10_ipd)

   begin
    if (REN_ipd = '1' ) then
	RD_ADD(4) <= RAD14_ipd;
	RD_ADD(3) <= RAD13_ipd;
	RD_ADD(2) <= RAD12_ipd;
	RD_ADD(1) <= RAD11_ipd;
	RD_ADD(0) <= RAD10_ipd;
    else
	RD_ADD <= x_add;
    end if;

    if (REN_ipd = '1' ) then
	RD_ADD2(4) <= RAD24_ipd;
	RD_ADD2(3) <= RAD23_ipd;
	RD_ADD2(2) <= RAD22_ipd;
	RD_ADD2(1) <= RAD21_ipd;
	RD_ADD2(0) <= RAD20_ipd;
    else
	RD_ADD2 <= x_add;
    end if;

   end process;


  VITALBehavior : PROCESS ( REN_ipd, OE_ipd, RAD24_ipd, RAD23_ipd, RAD22_ipd, RAD21_ipd, RAD20_ipd, RAD14_ipd, RAD13_ipd, RAD12_ipd, RAD11_ipd, RAD10_ipd)


   -- Temporary variables
   VARIABLE tmp_data : std_logic_vector (3 downto 0);
   VARIABLE readdata : LINE;
   VARIABLE first : boolean := TRUE;
   VARIABLE rd_address 		: integer := 0;
   VARIABLE rd_address_w 	: integer := 0;
   VARIABLE rd1 	: std_logic_vector(4 downto 0) ;
   VARIABLE rd2 	: std_logic_vector(4 downto 0) ;
   VARIABLE T 	: integer := 0;
   VARIABLE rd_viol_flag 	: X01 := '0';
   VARIABLE rd_viol_flag_w 	: X01 := '0';

    -------------------------------------------------------------------
    -- Functionality Section
    -------------------------------------------------------------------

BEGIN
if (first) then
          while( not(endfile(STF)) ) loop
                readline(STF,readdata) ;
                read(readdata,tmp_data) ;

    memory_array(T) <= tmp_data;
   T := T + 1;
  end loop;
end if;



rd1(4) := RAD14_ipd;
rd1(3) := RAD13_ipd;
rd1(2) := RAD12_ipd;
rd1(1) := RAD11_ipd;
rd1(0) := RAD10_ipd;
rd2(4) := RAD24_ipd;
rd2(3) := RAD23_ipd;
rd2(2) := RAD22_ipd;
rd2(1) := RAD21_ipd;
rd2(0) := RAD20_ipd;
-- READ CYCLE VIOLATION EFFECT

    if((RAD14_ipd'EVENT or RAD13_ipd'EVENT or RAD12_ipd'EVENT or RAD11_ipd'EVENT or RAD10_ipd'EVENT)  and REN_ipd = '1' and vecX(rd1)) then
	data_out <= x_data;
    elsif

-- VALID MEMORY READ


     ((RAD14_ipd'EVENT or RAD13_ipd'EVENT or RAD12_ipd'EVENT or RAD11_ipd'EVENT or RAD10_ipd'EVENT) and REN_ipd = '1' and not (vecX(rd1))) then
	rd_address := vec2int(rd1);
	data_out <= TRANSPORT memory_array(rd_address) ;
    end if;



    if((RAD24_ipd'EVENT or RAD23_ipd'EVENT or RAD22_ipd'EVENT or RAD21_ipd'EVENT or RAD20_ipd'EVENT)  and REN_ipd = '1' and vecX(rd2)) then
        data_out_w <= x_data;
    elsif

-- VALID MEMORY READ

     ((((RAD24_ipd'EVENT or RAD23_ipd'EVENT or RAD22_ipd'EVENT or RAD21_ipd'EVENT or RAD20_ipd'EVENT) and OE_ipd = '1' ) or ( OE_ipd = '1' and OE_ipd'EVENT )) and REN_ipd = '1' and not(rd_viol_flag_w = 'X') and not(vecX(rd2))) then
	rd_address_w := vec2int(rd2);
	data_out_w <= TRANSPORT memory_array(rd_address_w);
    end if;


  END PROCESS;

    -------------------------------------------------------------------------------
    -- Temporary output signal should get assigned to the output signal.
    -------------------------------------------------------------------------------


  PROCESS(data_out, RAD14_ipd, RAD13_ipd, RAD12_ipd, RAD11_ipd, RAD10_ipd)

     VARIABLE RDATA10_1 : std_logic := 'X';
     VARIABLE RDATA11_1 : std_logic := 'X';
     VARIABLE RDATA12_1 : std_logic := 'X';
     VARIABLE RDATA13_1 : std_logic := 'X';
     VARIABLE GLITCH1 : VitalGlitchDataType ;
    BEGIN
     RDATA10_1 := VitalBUF(data_out(0));
     RDATA11_1 := VitalBUF(data_out(1));
     RDATA12_1 := VitalBUF(data_out(2));
     RDATA13_1 := VitalBUF(data_out(3));

     VitalPathDelay01 ( RDATA13, GLITCH1, "RDATA13", RDATA13_1,
        Paths => (
        0 => ( RAD14_ipd'LAST_EVENT, tpd_RAD14_RDATA13, TRUE ),
        1 => ( RAD13_ipd'LAST_EVENT, tpd_RAD13_RDATA13, TRUE ),
        2 => ( RAD12_ipd'LAST_EVENT, tpd_RAD12_RDATA13, TRUE ),
        3 => ( RAD11_ipd'LAST_EVENT, tpd_RAD11_RDATA13, TRUE ),
        4 => ( RAD10_ipd'LAST_EVENT, tpd_RAD10_RDATA13, TRUE )),
        DefaultDelay=>VitalZeroDelay01,
        Mode=>VitalInertial,
        XON=>TRUE,
        MsgOn=>TRUE,
        MsgSeverity=>WARNING );

     VitalPathDelay01 ( RDATA12, GLITCH1, "RDATA12", RDATA12_1,
        Paths => (
        0 => ( RAD14_ipd'LAST_EVENT, tpd_RAD14_RDATA12, TRUE ),
        1 => ( RAD13_ipd'LAST_EVENT, tpd_RAD13_RDATA12, TRUE ),
        2 => ( RAD12_ipd'LAST_EVENT, tpd_RAD12_RDATA12, TRUE ),
        3 => ( RAD11_ipd'LAST_EVENT, tpd_RAD11_RDATA12, TRUE ),
        4 => ( RAD10_ipd'LAST_EVENT, tpd_RAD10_RDATA12, TRUE )),
        DefaultDelay=>VitalZeroDelay01,
        Mode=>VitalInertial,
        XON=>TRUE,
        MsgOn=>TRUE,
        MsgSeverity=>WARNING );

     VitalPathDelay01 ( RDATA11, GLITCH1, "RDATA11", RDATA11_1,
        Paths => (
        0 => ( RAD14_ipd'LAST_EVENT, tpd_RAD14_RDATA11, TRUE ),
        1 => ( RAD13_ipd'LAST_EVENT, tpd_RAD13_RDATA11, TRUE ),
        2 => ( RAD12_ipd'LAST_EVENT, tpd_RAD12_RDATA11, TRUE ),
        3 => ( RAD11_ipd'LAST_EVENT, tpd_RAD11_RDATA11, TRUE ),
        4 => ( RAD10_ipd'LAST_EVENT, tpd_RAD10_RDATA11, TRUE )),
        DefaultDelay=>VitalZeroDelay01,
        Mode=>VitalInertial,
        XON=>TRUE,
        MsgOn=>TRUE,
        MsgSeverity=>WARNING );

     VitalPathDelay01 ( RDATA10, GLITCH1, "RDATA10", RDATA10_1,
        Paths => (
        0 => ( RAD14_ipd'LAST_EVENT, tpd_RAD14_RDATA10, TRUE ),
        1 => ( RAD13_ipd'LAST_EVENT, tpd_RAD13_RDATA10, TRUE ),
        2 => ( RAD12_ipd'LAST_EVENT, tpd_RAD12_RDATA10, TRUE ),
        3 => ( RAD11_ipd'LAST_EVENT, tpd_RAD11_RDATA10, TRUE ),
        4 => ( RAD10_ipd'LAST_EVENT, tpd_RAD10_RDATA10, TRUE )),
        DefaultDelay=>VitalZeroDelay01,
        Mode=>VitalInertial,
        XON=>TRUE,
        MsgOn=>TRUE,
        MsgSeverity=>WARNING );

    END PROCESS;

  PROCESS(data_out_w, OE_ipd, RAD24_ipd, RAD23_ipd, RAD22_ipd, RAD21_ipd, RAD20_ipd)

     VARIABLE RDATA20_1 : std_logic := 'X';
     VARIABLE RDATA21_1 : std_logic := 'X';
     VARIABLE RDATA22_1 : std_logic := 'X';
     VARIABLE RDATA23_1 : std_logic := 'X';
     VARIABLE GLITCH2 : VitalGlitchDataType ;
    BEGIN
     RDATA20_1 := VitalBUF(data_out_w(0));
     RDATA21_1 := VitalBUF(data_out_w(1));
     RDATA22_1 := VitalBUF(data_out_w(2));
     RDATA23_1 := VitalBUF(data_out_w(3));

     VitalPathDelay01 ( RDATA23, GLITCH2, "RDATA23", RDATA23_1,
        Paths => (
        0 => ( RAD24_ipd'LAST_EVENT, tpd_RAD24_RDATA23, TRUE ),
        1 => ( RAD23_ipd'LAST_EVENT, tpd_RAD23_RDATA23, TRUE ),
        2 => ( RAD22_ipd'LAST_EVENT, tpd_RAD22_RDATA23, TRUE ),
        3 => ( RAD21_ipd'LAST_EVENT, tpd_RAD21_RDATA23, TRUE ),
        4 => ( RAD20_ipd'LAST_EVENT, tpd_RAD20_RDATA23, TRUE ),
        5 => ( OE_ipd'LAST_EVENT, tpd_OE_RDATA23, TRUE)),
        DefaultDelay=>VitalZeroDelay01,
        Mode=>VitalInertial,
        XON=>TRUE,
        MsgOn=>TRUE,
        MsgSeverity=>WARNING );

     VitalPathDelay01 ( RDATA22, GLITCH2, "RDATA22", RDATA22_1,
        Paths => (
        0 => ( RAD24_ipd'LAST_EVENT, tpd_RAD24_RDATA22, TRUE ),
        1 => ( RAD23_ipd'LAST_EVENT, tpd_RAD23_RDATA22, TRUE ),
        2 => ( RAD22_ipd'LAST_EVENT, tpd_RAD22_RDATA22, TRUE ),
        3 => ( RAD21_ipd'LAST_EVENT, tpd_RAD21_RDATA22, TRUE ),
        4 => ( RAD20_ipd'LAST_EVENT, tpd_RAD20_RDATA22, TRUE ),
        5 => ( OE_ipd'LAST_EVENT, tpd_OE_RDATA22, TRUE)),
        DefaultDelay=>VitalZeroDelay01,
        Mode=>VitalInertial,
        XON=>TRUE,
        MsgOn=>TRUE,
        MsgSeverity=>WARNING );

     VitalPathDelay01 ( RDATA21, GLITCH2, "RDATA21", RDATA21_1,
        Paths => (
        0 => ( RAD24_ipd'LAST_EVENT, tpd_RAD24_RDATA21, TRUE ),
        1 => ( RAD23_ipd'LAST_EVENT, tpd_RAD23_RDATA21, TRUE ),
        2 => ( RAD22_ipd'LAST_EVENT, tpd_RAD22_RDATA21, TRUE ),
        3 => ( RAD21_ipd'LAST_EVENT, tpd_RAD21_RDATA21, TRUE ),
        4 => ( RAD20_ipd'LAST_EVENT, tpd_RAD20_RDATA21, TRUE ),
        5 => ( OE_ipd'LAST_EVENT, tpd_OE_RDATA21, TRUE)),
        DefaultDelay=>VitalZeroDelay01,
        Mode=>VitalInertial,
        XON=>TRUE,
        MsgOn=>TRUE,
        MsgSeverity=>WARNING );

     VitalPathDelay01 ( RDATA20, GLITCH2, "RDATA20", RDATA20_1,
        Paths => (
        0 => ( RAD24_ipd'LAST_EVENT, tpd_RAD24_RDATA20, TRUE ),
        1 => ( RAD23_ipd'LAST_EVENT, tpd_RAD23_RDATA20, TRUE ),
        2 => ( RAD22_ipd'LAST_EVENT, tpd_RAD22_RDATA20, TRUE ),
        3 => ( RAD21_ipd'LAST_EVENT, tpd_RAD21_RDATA20, TRUE ),
        4 => ( RAD20_ipd'LAST_EVENT, tpd_RAD20_RDATA20, TRUE ),
        5 => ( OE_ipd'LAST_EVENT, tpd_OE_RDATA20, TRUE)),
        DefaultDelay=>VitalZeroDelay01,
        Mode=>VitalInertial,
        XON=>TRUE,
        MsgOn=>TRUE,
        MsgSeverity=>WARNING );

END PROCESS;


END VITAL_VF;
configuration CFG_R_DA_VITAL of R_DA is
        for VITAL_VF
        end for;
end CFG_R_DA_VITAL; 
-----------------------------------------------------------------------
-- VITAL model for R_DS 30.10 technology
-----------------------------------------------------------------------

LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.VITAL_timing.all;
USE IEEE.VITAL_primitives.all;
USE IEEE.std_logic_textio.all;
LIBRARY std;
USE std.textio.all;
LIBRARY VF1;
USE VF1.ALL;
USE VF1.RAMPACK.ALL;

-----------------------------------------------------------------------
-- ENTITY declaration
-----------------------------------------------------------------------

ENTITY R_DS IS
  GENERIC (
	tipd_REN		: VitalDelayType01			:= (0.0 ns, 0.0 ns);
	tipd_RCLK1		: VitalDelayType01			:= (0.0 ns, 0.0 ns);
	tipd_RCLK2		: VitalDelayType01			:= (0.0 ns, 0.0 ns);
	tipd_OE		: VitalDelayType01			:= (0.0 ns, 0.0 ns);
	tipd_RAD10		: VitalDelayType01	:= (0.0 ns, 0.0 ns);
	tipd_RAD11		: VitalDelayType01	:= (0.0 ns, 0.0 ns);
	tipd_RAD12		: VitalDelayType01	:= (0.0 ns, 0.0 ns);
	tipd_RAD13		: VitalDelayType01	:= (0.0 ns, 0.0 ns);
	tipd_RAD14		: VitalDelayType01	:= (0.0 ns, 0.0 ns);

	tipd_RAD20		: VitalDelayType01	:= (0.0 ns, 0.0 ns);
	tipd_RAD21		: VitalDelayType01	:= (0.0 ns, 0.0 ns);
	tipd_RAD22		: VitalDelayType01	:= (0.0 ns, 0.0 ns);
	tipd_RAD23		: VitalDelayType01	:= (0.0 ns, 0.0 ns);
	tipd_RAD24		: VitalDelayType01	:= (0.0 ns, 0.0 ns);

	tsetup_RAD10_RCLK1_noedge_posedge			: VitalDelayType := 1 ns;
	tsetup_RAD11_RCLK1_noedge_posedge			: VitalDelayType := 1 ns;
	tsetup_RAD12_RCLK1_noedge_posedge			: VitalDelayType := 1 ns;
	tsetup_RAD13_RCLK1_noedge_posedge			: VitalDelayType := 1 ns;
	tsetup_RAD14_RCLK1_noedge_posedge			: VitalDelayType := 1 ns;



	thold_RAD10_RCLK1_noedge_posedge			: VitalDelayType := 1 ns;
	thold_RAD11_RCLK1_noedge_posedge			: VitalDelayType := 1 ns;
	thold_RAD12_RCLK1_noedge_posedge			: VitalDelayType := 1 ns;
	thold_RAD13_RCLK1_noedge_posedge			: VitalDelayType := 1 ns;
	thold_RAD14_RCLK1_noedge_posedge			: VitalDelayType := 1 ns;


	tsetup_RAD20_RCLK2_noedge_posedge			: VitalDelayType := 1 ns;
	tsetup_RAD21_RCLK2_noedge_posedge			: VitalDelayType := 1 ns;
	tsetup_RAD22_RCLK2_noedge_posedge			: VitalDelayType := 1 ns;
	tsetup_RAD23_RCLK2_noedge_posedge			: VitalDelayType := 1 ns;
	tsetup_RAD24_RCLK2_noedge_posedge			: VitalDelayType := 1 ns;


	thold_RAD20_RCLK2_noedge_posedge			: VitalDelayType := 1 ns;
	thold_RAD21_RCLK2_noedge_posedge			: VitalDelayType := 1 ns;
	thold_RAD22_RCLK2_noedge_posedge			: VitalDelayType := 1 ns;
	thold_RAD23_RCLK2_noedge_posedge			: VitalDelayType := 1 ns;
	thold_RAD24_RCLK2_noedge_posedge			: VitalDelayType := 1 ns;

	tpd_RCLK1_RDATA10            			: VitalDelayType01 := (2 ns, 2 ns);
	tpd_RCLK1_RDATA11				: VitalDelayType01 := (2 ns, 2 ns);
	tpd_RCLK1_RDATA12				: VitalDelayType01 := (2 ns, 2 ns);
	tpd_RCLK1_RDATA13				: VitalDelayType01 := (2 ns, 2 ns);

	tpd_RCLK2_RDATA20				: VitalDelayType01 := (2 ns, 2 ns);
	tpd_RCLK2_RDATA21				: VitalDelayType01 := (2 ns, 2 ns);
	tpd_RCLK2_RDATA22				: VitalDelayType01 := (2 ns, 2 ns);
	tpd_RCLK2_RDATA23				: VitalDelayType01 := (2 ns, 2 ns);

	tpd_OE_RDATA20				: VitalDelayType01 := (2 ns, 2 ns);
	tpd_OE_RDATA21				: VitalDelayType01 := (2 ns, 2 ns);
	tpd_OE_RDATA22				: VitalDelayType01 := (2 ns, 2 ns);
	tpd_OE_RDATA23				: VitalDelayType01 := (2 ns, 2 ns);

	tpw_RCLK1_posedge					: VitalDelayType			:= 1 ns;
	tpw_RCLK2_posedge					: VitalDelayType			:= 1 ns;

	tsetup_REN_RCLK1_noedge_posedge			: VitalDelayType			:= 1 ns;
	tsetup_REN_RCLK2_noedge_posedge			: VitalDelayType			:= 1 ns;
	thold_REN_RCLK1_noedge_posedge			: VitalDelayType			:= 1 ns;
	thold_REN_RCLK2_noedge_posedge			: VitalDelayType			:= 1 ns;

	TimingChecksOn : BOOLEAN := TRUE;
	InstancePath : STRING := "*"
            );
  PORT	(
	REN		: IN	std_logic ;
	RCLK1		: IN	std_logic ;
	RCLK2		: IN	std_logic ;
	OE		: IN	std_logic ;
	RDATA20	        : OUT	std_logic := 'X';
	RDATA21	        : OUT	std_logic := 'X';
	RDATA22	        : OUT	std_logic := 'X';
	RDATA23	        : OUT	std_logic := 'X';
	RDATA10		: OUT	std_logic := 'X';
	RDATA11		: OUT	std_logic := 'X';
	RDATA12		: OUT	std_logic := 'X';
	RDATA13		: OUT	std_logic := 'X';
	RAD10		: IN	std_logic;
	RAD11		: IN	std_logic;
	RAD12		: IN	std_logic;
	RAD13		: IN	std_logic;
	RAD14		: IN	std_logic;
	RAD20		: IN	std_logic;
	RAD21		: IN	std_logic;
	RAD22		: IN	std_logic;
	RAD23		: IN	std_logic;
	RAD24		: IN	std_logic
	);


   ATTRIBUTE VITAL_LEVEL0 OF R_DS : ENTITY IS TRUE;

END R_DS;

-----------------------------------------------------------------------
-- ARCHITECTURE declaration
-----------------------------------------------------------------------
ARCHITECTURE VITAL_VF OF R_DS IS

    ATTRIBUTE VITAL_LEVEL1 OF VITAL_VF : ARCHITECTURE IS FALSE;

	file STF : text is in "rom_data";
	SIGNAL REN_ipd		: std_logic := 'X';
	SIGNAL RCLK1_ipd	: std_logic := '0';
	SIGNAL RCLK2_ipd	: std_logic := '0';
	SIGNAL RD_CLK		: std_logic := '0';
	SIGNAL RD_CLK_W		: std_logic := '0';
	SIGNAL OE_ipd	        : std_logic := 'X';
	SIGNAL RAD10_ipd	: std_logic;
	SIGNAL RAD11_ipd	: std_logic;
	SIGNAL RAD12_ipd	: std_logic;
	SIGNAL RAD13_ipd	: std_logic;
	SIGNAL RAD14_ipd	: std_logic;
	SIGNAL RD_ADD		: std_logic_vector(4 DOWNTO 0);
	SIGNAL RD_ADD_W		: std_logic_vector(4 DOWNTO 0);
	SIGNAL RAD20_ipd		: std_logic;
	SIGNAL RAD21_ipd		: std_logic;
	SIGNAL RAD22_ipd		: std_logic;
	SIGNAL RAD23_ipd		: std_logic;
	SIGNAL RAD24_ipd		: std_logic;
	SIGNAL data_out		: std_logic_vector(3 DOWNTO 0) := x_data;
	SIGNAL data_out_w	: std_logic_vector(3 DOWNTO 0) := x_data;
	SIGNAL output_delay_w	: time		:= 0 ns;
	SIGNAL output_delay	: time		:= 0 ns;

BEGIN
   
  ---------------------------------------------------------------------
  -- INPUT PATH DELAYs
  ---------------------------------------------------------------------
  WIREDELAY : BLOCK
  BEGIN
	VitalWireDelay (REN_ipd,		REN,		tipd_REN);
	VitalWireDelay (RCLK1_ipd,		RCLK1,		tipd_RCLK1);
	VitalWireDelay (RCLK2_ipd,		RCLK2,		tipd_RCLK2);
	VitalWireDelay (OE_ipd,			OE,		tipd_OE);
	VitalWireDelay (RAD10_ipd,		RAD10,		tipd_RAD10);
	VitalWireDelay (RAD11_ipd,		RAD11,		tipd_RAD11);
	VitalWireDelay (RAD12_ipd,		RAD12,		tipd_RAD12);
	VitalWireDelay (RAD13_ipd,		RAD13,		tipd_RAD13);
	VitalWireDelay (RAD14_ipd,		RAD14,		tipd_RAD14);
	VitalWireDelay (RAD20_ipd,		RAD20,		tipd_RAD20);
	VitalWireDelay (RAD21_ipd,		RAD21,		tipd_RAD21);
	VitalWireDelay (RAD22_ipd,		RAD22,		tipd_RAD22);
	VitalWireDelay (RAD23_ipd,		RAD23,		tipd_RAD23);
	VitalWireDelay (RAD24_ipd,		RAD24,		tipd_RAD24);

  END BLOCK;

  ---------------------------------------------------------------------
  -- Behavior Section
  ---------------------------------------------------------------------

  ---------------------------------------------------------------------
  -- Wrapper Section
  ---------------------------------------------------------------------

   wrapper_read_add : process(REN_ipd, OE_ipd, RAD10_ipd, RAD11_ipd, RAD12_ipd, RAD13_ipd, RAD14_ipd)

   begin
    if (REN_ipd = '1' ) then
	RD_ADD(0) <= RAD10_ipd;
	RD_ADD(1) <= RAD11_ipd;
	RD_ADD(2) <= RAD12_ipd;
	RD_ADD(3) <= RAD13_ipd;
	RD_ADD(4) <= RAD14_ipd;
    else
	RD_ADD <= x_add;
    end if;

   end process;

   wrapper_read_add_w : process(REN_ipd, OE_ipd, RAD20_ipd, RAD21_ipd, RAD22_ipd, RAD23_ipd, RAD24_ipd)

   begin
    if (REN_ipd = '1' ) then
	RD_ADD_W(0) <= RAD20_ipd;
	RD_ADD_W(1) <= RAD21_ipd;
	RD_ADD_W(2) <= RAD22_ipd;
	RD_ADD_W(3) <= RAD23_ipd;
	RD_ADD_W(4) <= RAD24_ipd;
    else
	RD_ADD_W <= x_add;
    end if;

   end process;

   wrapper_read_clk : process(REN_ipd, OE_ipd, RCLK1_ipd)

   begin
    if (REN_ipd = '1') then
	RD_CLK <= RCLK1_ipd;
    else
	RD_CLK <= '0';
    end if;

   end process;

   wrapper_read_clk_w : process(REN_ipd, OE_ipd, RCLK2_ipd)

   begin
    if (REN_ipd = '1' ) then
	RD_CLK_W <= RCLK2_ipd;
    else
	RD_CLK_W <= '0';
    end if;

   end process;


  VITALBehavior : PROCESS ( REN_ipd, RD_CLK_W, RD_CLK, RD_ADD, RD_ADD_W)

   VARIABLE memory_array : memory_array_typ;
--   VARIABLE array_data_out : data_word_typ := x_data;
--   VARIABLE array_data_out_w : data_word_typ := z_data;

   -- Temporary variables
   VARIABLE tmp_data : std_logic_vector (3 downto 0);
   VARIABLE readdata : LINE;
   VARIABLE first : boolean := TRUE;
   VARIABLE rd_address : integer := 0;
   VARIABLE T : integer := 0;
   VARIABLE rd_address_w : integer := 0;

   -- Timing Check results
   VARIABLE Pviol_RCLK				: std_logic := '0';
   VARIABLE PeriodData_RCLK			: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_RCLK_W			: std_logic := '0';
   VARIABLE PeriodData_RCLK_W			: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_RD_ADD_W_stp_hld_0		: std_logic := '0';
   VARIABLE TimingData_RD_ADD_W_stp_hld_0	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_RD_ADD_W_stp_hld_1		: std_logic := '0';
   VARIABLE TimingData_RD_ADD_W_stp_hld_1	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_RD_ADD_W_stp_hld_2		: std_logic := '0';
   VARIABLE TimingData_RD_ADD_W_stp_hld_2	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_RD_ADD_W_stp_hld_3		: std_logic := '0';
   VARIABLE TimingData_RD_ADD_W_stp_hld_3	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_RD_ADD_W_stp_hld_4		: std_logic := '0';
   VARIABLE TimingData_RD_ADD_W_stp_hld_4	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_RD_ADD_stp_hld_0		: std_logic := '0';
   VARIABLE TimingData_RD_ADD_stp_hld_0		: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_RD_ADD_stp_hld_1		: std_logic := '0';
   VARIABLE TimingData_RD_ADD_stp_hld_1		: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_RD_ADD_stp_hld_2		: std_logic := '0';
   VARIABLE TimingData_RD_ADD_stp_hld_2		: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_RD_ADD_stp_hld_3		: std_logic := '0';
   VARIABLE TimingData_RD_ADD_stp_hld_3		: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_RD_ADD_stp_hld_4		: std_logic := '0';
   VARIABLE TimingData_RD_ADD_stp_hld_4		: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_REN_hld			: std_logic := '0';
   VARIABLE TimingData_REN_hld			: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_REN_W_hld			: std_logic := '0';
   VARIABLE TimingData_REN_W_hld		: VitalTimingDataType := VitalTimingDataInit;



 BEGIN
    -------------------------------------------------------------------
    -- Timing Check Section
    -------------------------------------------------------------------
    IF (TimingChecksOn) THEN

	VitalPeriodPulseCheck  (Pviol_RCLK,
				PeriodData_RCLK,
				RD_CLK, "RCLK1",
				0.0 ns,
				0.0 ns,
				tpw_RCLK1_posedge,
				0.0 ns,
				TRUE,
				InstancePath & "/R_DS",
				TRUE,
				TRUE,
				WARNING );

	VitalPeriodPulseCheck  (Pviol_RCLK_W,
				PeriodData_RCLK_W,
				RD_CLK_W, "RCLK2",
				0.0 ns,
				0.0 ns,
				tpw_RCLK2_posedge,
				0.0 ns,
				TRUE,
				InstancePath & "/R_DS",
				TRUE,
				TRUE,
				WARNING );

	VitalSetupHoldCheck    (Tviol_RD_ADD_stp_hld_0,
				TimingData_RD_ADD_stp_hld_0,
				RD_ADD(0), "RAD10",
				0.0 ns,
				RD_CLK, "RCLK1",
				0.0 ns,
				tsetup_RAD10_RCLK1_noedge_posedge, tsetup_RAD10_RCLK1_noedge_posedge, 
				thold_RAD10_RCLK1_noedge_posedge, thold_RAD10_RCLK1_noedge_posedge,
				REN_ipd = '1',
				'/',
				InstancePath & "/R_DS",
				TRUE,
				TRUE,
				WARNING );

	VitalSetupHoldCheck    (Tviol_RD_ADD_stp_hld_1,
				TimingData_RD_ADD_stp_hld_1,
				RD_ADD(1), "RAD11",
				0.0 ns,
				RD_CLK, "RCLK1",
				0.0 ns,
				tsetup_RAD11_RCLK1_noedge_posedge, tsetup_RAD11_RCLK1_noedge_posedge,
				thold_RAD11_RCLK1_noedge_posedge, thold_RAD11_RCLK1_noedge_posedge,
				REN_ipd = '1',
				'R',
				InstancePath & "/R_DS",
				TRUE,
				TRUE,
				WARNING );

	VitalSetupHoldCheck    (Tviol_RD_ADD_stp_hld_2,
				TimingData_RD_ADD_stp_hld_2,
				RD_ADD(2), "RAD12",
				0.0 ns,
				RD_CLK, "RCLK1",
				0.0 ns,
				tsetup_RAD12_RCLK1_noedge_posedge, tsetup_RAD12_RCLK1_noedge_posedge,
				thold_RAD12_RCLK1_noedge_posedge, thold_RAD12_RCLK1_noedge_posedge,
				REN_ipd = '1',
				'/',
				InstancePath & "/R_DS",
				TRUE,
				TRUE,
				WARNING );

	VitalSetupHoldCheck    (Tviol_RD_ADD_stp_hld_3,
				TimingData_RD_ADD_stp_hld_3,
				RD_ADD(3), "RAD13",
				0.0 ns,
				RD_CLK, "RCLK1",
				0.0 ns,
				tsetup_RAD13_RCLK1_noedge_posedge, tsetup_RAD13_RCLK1_noedge_posedge,
				thold_RAD13_RCLK1_noedge_posedge, thold_RAD13_RCLK1_noedge_posedge,
				REN_ipd = '1',
				'/',
				InstancePath & "/R_DS",
				TRUE,
				TRUE,
				WARNING );

	VitalSetupHoldCheck    (Tviol_RD_ADD_stp_hld_4,
				TimingData_RD_ADD_stp_hld_4,
				RD_ADD(4), "RAD14",
				0.0 ns,
				RD_CLK, "RCLK1",
				0.0 ns,
				tsetup_RAD14_RCLK1_noedge_posedge, tsetup_RAD14_RCLK1_noedge_posedge,
				thold_RAD14_RCLK1_noedge_posedge, thold_RAD14_RCLK1_noedge_posedge,
				REN_ipd = '1',
				'/',
				InstancePath & "/R_DS",
				TRUE,
				TRUE,
				WARNING );

	VitalSetupHoldCheck    (Tviol_RD_ADD_W_stp_hld_0,
				TimingData_RD_ADD_W_stp_hld_0,
				RD_ADD_W(0), "RAD20",
				0.0 ns,
				RD_CLK_W, "RCLK2",
				0.0 ns,
				tsetup_RAD20_RCLK2_noedge_posedge, tsetup_RAD20_RCLK2_noedge_posedge,
				thold_RAD20_RCLK2_noedge_posedge, thold_RAD20_RCLK2_noedge_posedge,
				REN_ipd = '1',
				'/',
				InstancePath & "/R_DS",
				TRUE,
				TRUE,
				WARNING );

	VitalSetupHoldCheck    (Tviol_RD_ADD_W_stp_hld_1,
				TimingData_RD_ADD_W_stp_hld_1,
				RD_ADD_W(1), "RAD21",
				0.0 ns,
				RD_CLK_W, "RCLK2",
				0.0 ns,
				tsetup_RAD21_RCLK2_noedge_posedge, tsetup_RAD21_RCLK2_noedge_posedge,
				thold_RAD21_RCLK2_noedge_posedge, thold_RAD21_RCLK2_noedge_posedge,
				REN_ipd = '1',
				'/',
				InstancePath & "/R_DS",
				TRUE,
				TRUE,
				WARNING );

	VitalSetupHoldCheck    (Tviol_RD_ADD_W_stp_hld_2,
				TimingData_RD_ADD_W_stp_hld_2,
				RD_ADD_W(2), "RAD22",
				0.0 ns,
				RD_CLK_W, "RCLK2",
				0.0 ns,
				tsetup_RAD22_RCLK2_noedge_posedge,tsetup_RAD22_RCLK2_noedge_posedge, 
				thold_RAD22_RCLK2_noedge_posedge, thold_RAD22_RCLK2_noedge_posedge,
				REN_ipd = '1',
				'/',
				InstancePath & "/R_DS",
				TRUE,
				TRUE,
				WARNING );

	VitalSetupHoldCheck    (Tviol_RD_ADD_W_stp_hld_3,
				TimingData_RD_ADD_W_stp_hld_3,
				RD_ADD_W(3), "RAD23",
				0.0 ns,
				RD_CLK_W, "RCLK2",
				0.0 ns,
				tsetup_RAD23_RCLK2_noedge_posedge, tsetup_RAD23_RCLK2_noedge_posedge,
				thold_RAD23_RCLK2_noedge_posedge, thold_RAD23_RCLK2_noedge_posedge,
				REN_ipd = '1',
				'/',
				InstancePath & "/R_DS",
				TRUE,
				TRUE,
				WARNING );

	VitalSetupHoldCheck    (Tviol_RD_ADD_W_stp_hld_4,
				TimingData_RD_ADD_W_stp_hld_4,
				RD_ADD_W(4), "RAD24",
				0.0 ns,
				RD_CLK_W, "RCLK2",
				0.0 ns,
				tsetup_RAD24_RCLK2_noedge_posedge, tsetup_RAD24_RCLK2_noedge_posedge,
				thold_RAD24_RCLK2_noedge_posedge, thold_RAD24_RCLK2_noedge_posedge,
				REN_ipd = '1',
				'/',
				InstancePath & "/R_DS",
				TRUE,
				TRUE,
				WARNING );

	VitalSetupHoldCheck    (Tviol_REN_hld,
				TimingData_REN_hld,
				REN_ipd, "REN",
				0.0 ns,
				RD_CLK, "RCLK1",
				0.0 ns,
				tsetup_REN_RCLK1_noedge_posedge, tsetup_REN_RCLK1_noedge_posedge,
				thold_REN_RCLK1_noedge_posedge, thold_REN_RCLK1_noedge_posedge,
				True,
				'/',
				InstancePath & "/R_DS",
				TRUE,
				TRUE,
				WARNING );

	VitalSetupHoldCheck    (Tviol_REN_W_hld,
				TimingData_REN_W_hld,
				REN_ipd, "REN",
				0.0 ns,
				RD_CLK_W, "RCLK2",
				0.0 ns,
				tsetup_REN_RCLK2_noedge_posedge, tsetup_REN_RCLK2_noedge_posedge,
				thold_REN_RCLK2_noedge_posedge, thold_REN_RCLK2_noedge_posedge,
				True,
				'/',
				InstancePath & "/R_DS",
				TRUE,
				TRUE,
				WARNING );

    END IF; -- Timing Check Section

    -------------------------------------------------------------------
    -- Functionality Section
    -------------------------------------------------------------------


if (first) then
          while( not(endfile(STF)) ) loop
                readline(STF,readdata) ;
                read(readdata,tmp_data) ;

--  for T in 0 to 31 loop
 --   READLINE (STF,readdata);
  --  Read (readdata,tmp_data);
    memory_array(T) := tmp_data;
   T := T + 1;
  end loop;
end if;


-- READ ADDRESS CYCLE VIOLATION EFFECT

    if( Tviol_RD_ADD_stp_hld_0 = 'X' or Tviol_RD_ADD_stp_hld_1 = 'X' or Tviol_RD_ADD_stp_hld_2 = 'X' or Tviol_RD_ADD_stp_hld_3 = 'X' or Tviol_RD_ADD_stp_hld_4 = 'X' or Pviol_RCLK = 'X' or Tviol_REN_hld = 'X' or (RD_CLK'EVENT and RD_CLK = '1' and vecX(RD_ADD))) then
	--output_delay <= 0 ns;
	data_out <= x_data;
    elsif


-- VALID MEMORY READ

    (RD_CLK'EVENT and RD_CLK = '1' and not( Tviol_RD_ADD_stp_hld_0 = 'X' or Tviol_RD_ADD_stp_hld_1 = 'X' or Tviol_RD_ADD_stp_hld_2 = 'X' or Tviol_RD_ADD_stp_hld_3 = 'X' or Tviol_RD_ADD_stp_hld_4 = 'X' or Pviol_RCLK = 'X' or Tviol_REN_hld = 'X' or vecX(RD_ADD) )) then
	rd_address := vec2int(RD_ADD);
	--output_delay <= tpd_RCLK1_RDATA1_posedge(0);
	data_out <= memory_array(rd_address);
    end if;

    if RD_CLK'EVENT and RD_CLK /= RCLK1_ipd and RD_CLK'LAST_VALUE = '1' then
	--output_delay <= 0 ns;
	data_out <= x_data;
    end if;


-- READ ADDRESS CYCLE VIOLATION EFFECT

    if( Tviol_RD_ADD_W_stp_hld_0 = 'X' or Tviol_RD_ADD_W_stp_hld_1 = 'X' or Tviol_RD_ADD_W_stp_hld_2 = 'X' or Tviol_RD_ADD_W_stp_hld_3 = 'X' or Tviol_RD_ADD_W_stp_hld_4 = 'X' or Pviol_RCLK_W = 'X' or Tviol_REN_W_hld = 'X' or (RD_CLK_W'EVENT and RD_CLK_W = '1' and vecX(RD_ADD_W)) ) then
	--output_delay_w <= 0 ns;
	data_out_w <= x_data;
    elsif

-- VALID MEMORY READ

    (RD_CLK_W'EVENT and RD_CLK_W = '1' and not( Tviol_RD_ADD_W_stp_hld_0 = 'X' or Tviol_RD_ADD_W_stp_hld_1 = 'X' or Tviol_RD_ADD_W_stp_hld_2 = 'X' or Tviol_RD_ADD_W_stp_hld_3 = 'X' or Tviol_RD_ADD_W_stp_hld_4 = 'X' or Pviol_RCLK_W = 'X' or Tviol_REN_W_hld = 'X' or vecX(RD_ADD_W) ))then
	rd_address_w := vec2int(RD_ADD_W);
	--output_delay_w <= tpd_RCLK2_RDATA2_posedge(0);
	data_out_w <= memory_array(rd_address_w);
    end if;

    if RD_CLK_W'EVENT and RD_CLK_W /= RCLK2_ipd and RD_CLK_W'LAST_VALUE = '1' then
	--output_delay_w <= 0 ns;
	data_out_w <= x_data;
    end if;

--data_out <= array_data_out;

--data_out_w <= array_data_out_w;


  END PROCESS;

    -------------------------------------------------------------------------------
    -- Temporary output signal should get assigned to the output signal.
    -------------------------------------------------------------------------------

  PROCESS(data_out, RCLK1_ipd)

     VARIABLE RDATA13_1 :std_logic := 'X';
     VARIABLE RDATA12_1 :std_logic := 'X';
     VARIABLE RDATA11_1 :std_logic := 'X';
     VARIABLE RDATA10_1 :std_logic := 'X';
     VARIABLE GLITCH1 : VitalGlitchDataType ;

    BEGIN

       RDATA13_1 := VitalBUF(data_out(3));
       RDATA12_1 := VitalBUF(data_out(2));
       RDATA11_1 := VitalBUF(data_out(1));
       RDATA10_1 := VitalBUF(data_out(0));

     VitalPathDelay01 ( RDATA13, GLITCH1, "RDATA13", RDATA13_1,
        Paths => (
        0 => ( RCLK1_ipd'LAST_EVENT, tpd_RCLK1_RDATA13, TRUE )),
        DefaultDelay=>VitalZeroDelay01,
        Mode=>VitalInertial,
        XON=>TRUE,
        MsgOn=>TRUE,
        MsgSeverity=>WARNING );

     VitalPathDelay01 ( RDATA12, GLITCH1, "RDATA12", RDATA12_1,
        Paths => (
        0 => ( RCLK1_ipd'LAST_EVENT, tpd_RCLK1_RDATA12, TRUE )),
        DefaultDelay=>VitalZeroDelay01,
        Mode=>VitalInertial,
        XON=>TRUE,
        MsgOn=>TRUE,
        MsgSeverity=>WARNING );

     VitalPathDelay01 ( RDATA11, GLITCH1, "RDATA11", RDATA11_1,
        Paths => (
        0 => ( RCLK1_ipd'LAST_EVENT, tpd_RCLK1_RDATA11, TRUE )),
        DefaultDelay=>VitalZeroDelay01,
        Mode=>VitalInertial,
        XON=>TRUE,
        MsgOn=>TRUE,
        MsgSeverity=>WARNING );

     VitalPathDelay01 ( RDATA10, GLITCH1, "RDATA10", RDATA10_1,
        Paths => (
        0 => ( RCLK1_ipd'LAST_EVENT, tpd_RCLK1_RDATA10, TRUE )),
        DefaultDelay=>VitalZeroDelay01,
        Mode=>VitalInertial,
        XON=>TRUE,
        MsgOn=>TRUE,
        MsgSeverity=>WARNING );


     
    END PROCESS;

  PROCESS(data_out_w, RCLK2_ipd, OE_ipd)

     VARIABLE RDATA23_1 :std_logic := 'X';
     VARIABLE RDATA22_1 :std_logic := 'X';
     VARIABLE RDATA21_1 :std_logic := 'X';
     VARIABLE RDATA20_1 :std_logic := 'X';
     VARIABLE GLITCH2 : VitalGlitchDataType ;

    BEGIN

       RDATA23_1 := VitalBUF(data_out_w(3));
       RDATA22_1 := VitalBUF(data_out_w(2));
       RDATA21_1 := VitalBUF(data_out_w(1));
       RDATA20_1 := VitalBUF(data_out_w(0));

     VitalPathDelay01 ( RDATA23, GLITCH2, "RDATA23", RDATA23_1,
        Paths => (
        0 => ( RCLK2_ipd'LAST_EVENT, tpd_RCLK2_RDATA23, TRUE ),
        1 => ( OE_ipd'LAST_EVENT, tpd_OE_RDATA23, TRUE)),
        DefaultDelay=>VitalZeroDelay01,
        Mode=>VitalInertial,
        XON=>TRUE,
        MsgOn=>TRUE,
        MsgSeverity=>WARNING );

     VitalPathDelay01 ( RDATA22, GLITCH2, "RDATA22", RDATA22_1,
        Paths => (
        0 => ( RCLK2_ipd'LAST_EVENT, tpd_RCLK2_RDATA22, TRUE ),
        1 => ( OE_ipd'LAST_EVENT, tpd_OE_RDATA22, TRUE)),
        DefaultDelay=>VitalZeroDelay01,
        Mode=>VitalInertial,
        XON=>TRUE,
        MsgOn=>TRUE,
        MsgSeverity=>WARNING );

     VitalPathDelay01 ( RDATA21, GLITCH2, "RDATA21", RDATA21_1,
        Paths => (
        0 => ( RCLK2_ipd'LAST_EVENT, tpd_RCLK2_RDATA21, TRUE ),
        1 => ( OE_ipd'LAST_EVENT, tpd_OE_RDATA21, TRUE)),
        DefaultDelay=>VitalZeroDelay01,
        Mode=>VitalInertial,
        XON=>TRUE,
        MsgOn=>TRUE,
        MsgSeverity=>WARNING );

     VitalPathDelay01 ( RDATA20, GLITCH2, "RDATA20", RDATA20_1,
        Paths => (
        0 => ( RCLK2_ipd'LAST_EVENT, tpd_RCLK2_RDATA20, TRUE ),
        1 => ( OE_ipd'LAST_EVENT, tpd_OE_RDATA20, TRUE)),
        DefaultDelay=>VitalZeroDelay01,
        Mode=>VitalInertial,
        XON=>TRUE,
        MsgOn=>TRUE,
        MsgSeverity=>WARNING );

END PROCESS;
     

END VITAL_VF;
configuration CFG_R_DS_VITAL of R_DS is
        for VITAL_VF
        end for;
end CFG_R_DS_VITAL;
-----------------------------------------------------------------------


-----------------------------------------------------------------------
-- VITAL model for R_SA 30.10 technology
-----------------------------------------------------------------------

LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.VITAL_timing.all;
USE IEEE.VITAL_primitives.all;
USE IEEE.std_logic_textio.all;
LIBRARY std;
USE std.textio.all;
LIBRARY VF1;
USE VF1.ALL;
USE VF1.RAMPACK.ALL;

-----------------------------------------------------------------------
-- ENTITY declaration
-----------------------------------------------------------------------

ENTITY R_SA IS
  GENERIC (
	tipd_REN		: VitalDelayType01	:= (0.0 ns, 0.0 ns);
	tipd_RAD0		: VitalDelayType01	:= (0.0 ns, 0.0 ns);
	tipd_RAD1		: VitalDelayType01	:= (0.0 ns, 0.0 ns);
	tipd_RAD2		: VitalDelayType01	:= (0.0 ns, 0.0 ns);
	tipd_RAD3		: VitalDelayType01	:= (0.0 ns, 0.0 ns);
	tipd_RAD4		: VitalDelayType01	:= (0.0 ns, 0.0 ns);


	tpd_RAD0_RDATA0					: VitalDelayType01 := (2 ns,2 ns);
	tpd_RAD0_RDATA1					: VitalDelayType01 := (2 ns,2 ns);
	tpd_RAD0_RDATA2					: VitalDelayType01 := (2 ns,2 ns);
	tpd_RAD0_RDATA3					: VitalDelayType01 := (2 ns,2 ns);
	tpd_RAD1_RDATA0					: VitalDelayType01 := (2 ns,2 ns);
	tpd_RAD1_RDATA1					: VitalDelayType01 := (2 ns,2 ns);
	tpd_RAD1_RDATA2					: VitalDelayType01 := (2 ns,2 ns);
	tpd_RAD1_RDATA3					: VitalDelayType01 := (2 ns,2 ns);
	tpd_RAD2_RDATA0					: VitalDelayType01 := (2 ns,2 ns);
	tpd_RAD2_RDATA1					: VitalDelayType01 := (2 ns,2 ns);
	tpd_RAD2_RDATA2					: VitalDelayType01 := (2 ns,2 ns);
	tpd_RAD2_RDATA3					: VitalDelayType01 := (2 ns,2 ns);
	tpd_RAD3_RDATA0					: VitalDelayType01 := (2 ns,2 ns);
	tpd_RAD3_RDATA1					: VitalDelayType01 := (2 ns,2 ns);
	tpd_RAD3_RDATA2					: VitalDelayType01 := (2 ns,2 ns);
	tpd_RAD3_RDATA3					: VitalDelayType01 := (2 ns,2 ns);
	tpd_RAD4_RDATA0					: VitalDelayType01 := (2 ns,2 ns);
	tpd_RAD4_RDATA1					: VitalDelayType01 := (2 ns,2 ns);
	tpd_RAD4_RDATA2					: VitalDelayType01 := (2 ns,2 ns);
	tpd_RAD4_RDATA3					: VitalDelayType01 := (2 ns,2 ns);

	tpd_REN_RDATA0					: VitalDelayType01 := (2 ns,2 ns);
	tpd_REN_RDATA1					: VitalDelayType01 := (2 ns,2 ns);
	tpd_REN_RDATA2					: VitalDelayType01 := (2 ns,2 ns);
	tpd_REN_RDATA3					: VitalDelayType01 := (2 ns,2 ns);
	TimingChecksOn : BOOLEAN := TRUE;
	InstancePath : STRING := "*"
            );
  PORT	(
	REN		: IN	std_logic ;
	RDATA0		: OUT	std_logic;
	RDATA1		: OUT	std_logic;
	RDATA2		: OUT	std_logic;
	RDATA3		: OUT	std_logic;

	RAD0		: IN	std_logic;
	RAD1		: IN	std_logic;
	RAD2		: IN	std_logic;
	RAD3		: IN	std_logic;
	RAD4		: IN	std_logic
	);


   ATTRIBUTE VITAL_LEVEL0 OF R_SA : ENTITY IS TRUE;

END R_SA;

-----------------------------------------------------------------------
-- ARCHITECTURE declaration
-----------------------------------------------------------------------
ARCHITECTURE VITAL_VF OF R_SA IS

    ATTRIBUTE VITAL_LEVEL1 OF VITAL_VF : ARCHITECTURE IS FALSE;

	file STF : text is in "rom_data";
	SIGNAL REN_ipd		: std_logic := 'X';
	SIGNAL RAD0_ipd		: std_logic;
	SIGNAL RAD1_ipd		: std_logic;
	SIGNAL RAD2_ipd		: std_logic;
	SIGNAL RAD3_ipd		: std_logic;
	SIGNAL RAD4_ipd		: std_logic;

	SIGNAL RD_ADD		: std_logic_vector(4 DOWNTO 0);
	SIGNAL data_out		: std_logic_vector(3 DOWNTO 0) := x_data;
	SIGNAL output_delay	: time		:= 0 ns;
	SIGNAL memory_array	: memory_array_typ;

BEGIN
   
  ---------------------------------------------------------------------
  -- INPUT PATH DELAYs
  ---------------------------------------------------------------------
  WIREDELAY : BLOCK
  BEGIN
	VitalWireDelay (REN_ipd,		REN,		tipd_REN);
	VitalWireDelay (RAD0_ipd,		RAD0,		tipd_RAD0);
	VitalWireDelay (RAD1_ipd,		RAD1,		tipd_RAD1);
	VitalWireDelay (RAD2_ipd,		RAD2,		tipd_RAD2);
	VitalWireDelay (RAD3_ipd,		RAD3,		tipd_RAD3);
	VitalWireDelay (RAD4_ipd,		RAD4,		tipd_RAD4);

  END BLOCK;

  ---------------------------------------------------------------------
  -- Behavior Section
  ---------------------------------------------------------------------

  ---------------------------------------------------------------------
  -- Wrapper Section
  ---------------------------------------------------------------------

   wrapper_read_add : process(REN_ipd, RAD0_ipd, RAD1_ipd, RAD2_ipd, RAD3_ipd, RAD4_ipd)

   begin
    if (REN_ipd = '1' ) then
	RD_ADD(0) <= RAD0_ipd;
	RD_ADD(1) <= RAD1_ipd;
	RD_ADD(2) <= RAD2_ipd;
	RD_ADD(3) <= RAD3_ipd;
	RD_ADD(4) <= RAD4_ipd;
    else
	RD_ADD <= x_add;
    end if;

   end process;


  VITALBehavior : PROCESS ( REN_ipd, RD_ADD,  RAD0_ipd,  RAD1_ipd,  RAD2_ipd,  RAD3_ipd,  RAD4_ipd )


   -- Temporary variables
   VARIABLE tmp_data : std_logic_vector (3 downto 0);
   VARIABLE readdata : LINE;
   VARIABLE first : boolean := TRUE;
   VARIABLE rd_address 		: integer := 0;
   VARIABLE T 		: integer := 0;
   VARIABLE rd_viol_flag 	: X01 := '0';


    -------------------------------------------------------------------
    -- Functionality Section
    -------------------------------------------------------------------

BEGIN

if (first) then
          while( not(endfile(STF)) ) loop
                readline(STF,readdata) ;
                read(readdata,tmp_data) ;

    memory_array(T) <= tmp_data;
    T := T + 1;
  end loop;
first := FALSE;
end if;


-- READ CYCLE VIOLATION EFFECT

    if(RD_ADD'EVENT and REN_ipd = '1' and vecX(RD_ADD)) then
	--output_delay <= 0 ns;
	data_out <=  x_data;
    elsif

-- VALID MEMORY READ

   (((RD_ADD'EVENT and REN_ipd = '1' ) or (REN_ipd'EVENT and REN_ipd = '1')) and not (vecX(RD_ADD))) then
	rd_address := vec2int(RD_ADD);
	data_out <=  memory_array(rd_address) ;
    end if;


  END PROCESS;

    -------------------------------------------------------------------------------
    -- Temporary output signal should get assigned to the output signal.
    -------------------------------------------------------------------------------
    PROCESS(data_out, REN_ipd, RAD4_ipd, RAD3_ipd, RAD2_ipd, RAD1_ipd, RAD0_ipd)

      VARIABLE GLITCH : VitalGlitchDataType;
      VARIABLE RDATA3_1 : std_logic := 'X';
      VARIABLE RDATA2_1 : std_logic := 'X';
      VARIABLE RDATA1_1 : std_logic := 'X';
      VARIABLE RDATA0_1 : std_logic := 'X';

   BEGIN
       RDATA3_1 := VitalBUF(data_out(3));
       RDATA2_1 := VitalBUF(data_out(2));
       RDATA1_1 := VitalBUF(data_out(1));
       RDATA0_1 := VitalBUF(data_out(0));

     VitalPathDelay01 ( RDATA3, GLITCH, "RDATA3", RDATA3_1,
        Paths => (
        0 => ( REN_ipd'LAST_EVENT, tpd_REN_RDATA3, TRUE ),
        1 => ( RAD4_ipd'LAST_EVENT, tpd_RAD4_RDATA3, TRUE ),
        2 => ( RAD3_ipd'LAST_EVENT, tpd_RAD3_RDATA3, TRUE ),
        3 => ( RAD2_ipd'LAST_EVENT, tpd_RAD2_RDATA3, TRUE ),
        4 => ( RAD1_ipd'LAST_EVENT, tpd_RAD1_RDATA3, TRUE ),
        5 => ( RAD0_ipd'LAST_EVENT, tpd_RAD0_RDATA3, TRUE )),
        DefaultDelay=>VitalZeroDelay01,
        Mode=>VitalInertial,
        XON=>TRUE,
        MsgOn=>TRUE,
        MsgSeverity=>WARNING );

     VitalPathDelay01 ( RDATA2, GLITCH, "RDATA2", RDATA2_1,
        Paths => (
        0 => ( REN_ipd'LAST_EVENT, tpd_REN_RDATA2, TRUE ),
        1 => ( RAD4_ipd'LAST_EVENT, tpd_RAD4_RDATA2, TRUE ),
        2 => ( RAD3_ipd'LAST_EVENT, tpd_RAD3_RDATA2, TRUE ),
        3 => ( RAD2_ipd'LAST_EVENT, tpd_RAD2_RDATA2, TRUE ),
        4 => ( RAD1_ipd'LAST_EVENT, tpd_RAD1_RDATA2, TRUE ),
        5 => ( RAD0_ipd'LAST_EVENT, tpd_RAD0_RDATA2, TRUE )),
        DefaultDelay=>VitalZeroDelay01,
        Mode=>VitalInertial,
        XON=>TRUE,
        MsgOn=>TRUE,
        MsgSeverity=>WARNING );

     VitalPathDelay01 ( RDATA1, GLITCH, "RDATA1", RDATA1_1,
        Paths => (
        0 => ( REN_ipd'LAST_EVENT, tpd_REN_RDATA1, TRUE ),
        1 => ( RAD4_ipd'LAST_EVENT, tpd_RAD4_RDATA1, TRUE ),
        2 => ( RAD3_ipd'LAST_EVENT, tpd_RAD3_RDATA1, TRUE ),
        3 => ( RAD2_ipd'LAST_EVENT, tpd_RAD2_RDATA1, TRUE ),
        4 => ( RAD1_ipd'LAST_EVENT, tpd_RAD1_RDATA1, TRUE ),
        5 => ( RAD0_ipd'LAST_EVENT, tpd_RAD0_RDATA1, TRUE )),
        DefaultDelay=>VitalZeroDelay01,
        Mode=>VitalInertial,
        XON=>TRUE,
        MsgOn=>TRUE,
        MsgSeverity=>WARNING );

     VitalPathDelay01 ( RDATA0, GLITCH, "RDATA0", RDATA0_1,
        Paths => (
        0 => ( REN_ipd'LAST_EVENT, tpd_REN_RDATA0, TRUE ),
        1 => ( RAD4_ipd'LAST_EVENT, tpd_RAD4_RDATA0, TRUE ),
        2 => ( RAD3_ipd'LAST_EVENT, tpd_RAD3_RDATA0, TRUE ),
        3 => ( RAD2_ipd'LAST_EVENT, tpd_RAD2_RDATA0, TRUE ),
        4 => ( RAD1_ipd'LAST_EVENT, tpd_RAD1_RDATA0, TRUE ),
        5 => ( RAD0_ipd'LAST_EVENT, tpd_RAD0_RDATA0, TRUE )),
        DefaultDelay=>VitalZeroDelay01,
        Mode=>VitalInertial,
        XON=>TRUE,
        MsgOn=>TRUE,
        MsgSeverity=>WARNING );

END PROCESS;

END VITAL_VF;
configuration CFG_R_SA_VITAL of R_SA is
        for VITAL_VF
        end for;
end CFG_R_SA_VITAL;
-----------------------------------------------------------------------

-----------------------------------------------------------------------
-- VITAL model for R_SS 30.10 technology
-----------------------------------------------------------------------

LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.VITAL_timing.all;
USE IEEE.VITAL_primitives.all;
USE IEEE.std_logic_textio.all;
LIBRARY std;
USE std.textio.all;
LIBRARY VF1;
USE VF1.ALL;
USE VF1.RAMPACK.ALL;

-----------------------------------------------------------------------
-- ENTITY declaration
-----------------------------------------------------------------------

ENTITY R_SS IS
  GENERIC (
	tipd_REN		: VitalDelayType01			:= (0.0 ns, 0.0 ns);
	tipd_RCLK		: VitalDelayType01			:= (0.0 ns, 0.0 ns);
	tipd_RAD0		: VitalDelayType01	:= (0.0 ns, 0.0 ns);
	tipd_RAD1		: VitalDelayType01	:= (0.0 ns, 0.0 ns);
	tipd_RAD2		: VitalDelayType01	:= (0.0 ns, 0.0 ns);
	tipd_RAD3		: VitalDelayType01	:= (0.0 ns, 0.0 ns);
	tipd_RAD4		: VitalDelayType01	:= (0.0 ns, 0.0 ns);

	tsetup_RAD0_RCLK_noedge_posedge			: VitalDelayType := 1 ns;
	tsetup_RAD1_RCLK_noedge_posedge			: VitalDelayType := 1 ns;
	tsetup_RAD2_RCLK_noedge_posedge			: VitalDelayType := 1 ns;
	tsetup_RAD3_RCLK_noedge_posedge			: VitalDelayType := 1 ns;
	tsetup_RAD4_RCLK_noedge_posedge			: VitalDelayType := 1 ns;


	thold_RAD0_RCLK_noedge_posedge			: VitalDelayType := 1 ns;
	thold_RAD1_RCLK_noedge_posedge			: VitalDelayType := 1 ns;
	thold_RAD2_RCLK_noedge_posedge			: VitalDelayType := 1 ns;
	thold_RAD3_RCLK_noedge_posedge			: VitalDelayType := 1 ns;
	thold_RAD4_RCLK_noedge_posedge			: VitalDelayType := 1 ns;


	tpd_RCLK_RDATA0			: VitalDelayType01 := (2 ns,2 ns);
	tpd_RCLK_RDATA1			: VitalDelayType01 := (2 ns,2 ns);
	tpd_RCLK_RDATA2			: VitalDelayType01 := (2 ns,2 ns);
	tpd_RCLK_RDATA3			: VitalDelayType01 := (2 ns,2 ns);

	tpw_RCLK_posedge					: VitalDelayType			:= 1 ns;
	tsetup_REN_RCLK_noedge_posedge			: VitalDelayType			:= 1 ns;
	thold_REN_RCLK_noedge_posedge			: VitalDelayType			:= 1 ns;

	TimingChecksOn : BOOLEAN := TRUE;
	InstancePath : STRING := "*"
            );
  PORT	(
	REN		: IN	std_logic ;
	RCLK		: IN	std_logic ;
	RDATA0		: OUT	std_logic;
	RDATA1		: OUT	std_logic;
	RDATA2		: OUT	std_logic;
	RDATA3		: OUT	std_logic;
	RAD0		: IN	std_logic;
	RAD1		: IN	std_logic;
	RAD2		: IN	std_logic;
	RAD3		: IN	std_logic;
	RAD4		: IN	std_logic
	);


   ATTRIBUTE VITAL_LEVEL0 OF R_SS : ENTITY IS TRUE;

END R_SS;

-----------------------------------------------------------------------
-- ARCHITECTURE declaration
-----------------------------------------------------------------------
ARCHITECTURE VITAL_VF OF R_SS IS

    ATTRIBUTE VITAL_LEVEL1 OF VITAL_VF : ARCHITECTURE IS FALSE;

	file STF : text is in "rom_data";
	SIGNAL REN_ipd		: std_logic := 'X';
	SIGNAL RCLK_ipd		: std_logic := '0';
	SIGNAL RD_CLK		: std_logic := '0';
	SIGNAL RAD0_ipd		: std_logic;
	SIGNAL RAD1_ipd		: std_logic;
	SIGNAL RAD2_ipd		: std_logic;
	SIGNAL RAD3_ipd		: std_logic;
	SIGNAL RAD4_ipd		: std_logic;
	SIGNAL RD_ADD		: std_logic_vector(4 DOWNTO 0);
	SIGNAL data_out		: std_logic_vector(3 DOWNTO 0);
	SIGNAL output_delay	: time		:= 0 ns;

BEGIN
   
  ---------------------------------------------------------------------
  -- INPUT PATH DELAYs
  ---------------------------------------------------------------------
  WIREDELAY : BLOCK
  BEGIN
	VitalWireDelay (REN_ipd,		REN,		tipd_REN);
	VitalWireDelay (RCLK_ipd,		RCLK,		tipd_RCLK);
	VitalWireDelay (RAD0_ipd,		RAD0,		tipd_RAD0);
	VitalWireDelay (RAD1_ipd,		RAD1,		tipd_RAD1);
	VitalWireDelay (RAD2_ipd,		RAD2,		tipd_RAD2);
	VitalWireDelay (RAD3_ipd,		RAD3,		tipd_RAD3);
	VitalWireDelay (RAD4_ipd,		RAD4,		tipd_RAD4);

  END BLOCK;

  ---------------------------------------------------------------------
  -- Behavior Section
  ---------------------------------------------------------------------

  ---------------------------------------------------------------------
  -- Wrapper Section
  ---------------------------------------------------------------------

   wrapper_read_add : process(REN_ipd, RAD4_ipd, RAD3_ipd, RAD2_ipd, RAD1_ipd, RAD0_ipd)

   begin
    if (REN_ipd = '1' ) then
	RD_ADD(4) <= RAD4_ipd;
	RD_ADD(3) <= RAD3_ipd;
	RD_ADD(2) <= RAD2_ipd;
	RD_ADD(1) <= RAD1_ipd;
	RD_ADD(0) <= RAD0_ipd;
    else
	RD_ADD <= x_add;
    end if;

   end process;

   wrapper_read_clk : process(REN_ipd, RCLK_ipd)

   begin
    if (REN_ipd = '1' ) then
	RD_CLK <= RCLK_ipd;
    else
	RD_CLK <= '0';
    end if;

   end process;


  VITALBehavior : PROCESS ( REN_ipd, RD_CLK, RD_ADD)

   VARIABLE memory_array : memory_array_typ := (others =>(others=>'X'));

   -- Temporary variables
   VARIABLE tmp_data : std_logic_vector (3 downto 0);
   VARIABLE readdata : LINE;
   VARIABLE first : boolean := TRUE;
   VARIABLE rd_address : integer := 0;
   VARIABLE T : integer := 0;

   -- Timing Check results
   VARIABLE Pviol_RCLK			: std_logic := '0';
   VARIABLE PeriodData_RCLK		: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_RD_ADD_stp_hld_0	: std_logic := '0';
   VARIABLE TimingData_RD_ADD_stp_hld_0	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_RD_ADD_stp_hld_1	: std_logic := '0';
   VARIABLE TimingData_RD_ADD_stp_hld_1	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_RD_ADD_stp_hld_2	: std_logic := '0';
   VARIABLE TimingData_RD_ADD_stp_hld_2	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_RD_ADD_stp_hld_3	: std_logic := '0';
   VARIABLE TimingData_RD_ADD_stp_hld_3	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_RD_ADD_stp_hld_4	: std_logic := '0';
   VARIABLE TimingData_RD_ADD_stp_hld_4	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_REN_hld		: std_logic := '0';
   VARIABLE TimingData_REN_hld		: VitalTimingDataType := VitalTimingDataInit;



 BEGIN
    -------------------------------------------------------------------
    -- Timing Check Section
    -------------------------------------------------------------------
    IF (TimingChecksOn) THEN

	VitalPeriodPulseCheck  (Pviol_RCLK,
				PeriodData_RCLK,
				RD_CLK, "RCLK",
				0.0 ns,
				0.0 ns,
				tpw_RCLK_posedge,
				0.0 ns,
				REN_ipd = '1' ,
				InstancePath & "/R_SS",
				TRUE,
				TRUE,
				WARNING );

	VitalSetupHoldCheck    (Tviol_RD_ADD_stp_hld_0,
				TimingData_RD_ADD_stp_hld_0,
				RD_ADD(0), "RAD0",
				0.0 ns,
				RD_CLK, "RCLK",
				0.0 ns,
				tsetup_RAD0_RCLK_noedge_posedge, tsetup_RAD0_RCLK_noedge_posedge, 
				thold_RAD0_RCLK_noedge_posedge, thold_RAD0_RCLK_noedge_posedge,
				REN_ipd = '1' ,
				'/',
				InstancePath & "/R_SS",
				TRUE,
				TRUE,
				WARNING );

	VitalSetupHoldCheck    (Tviol_RD_ADD_stp_hld_1,
				TimingData_RD_ADD_stp_hld_1,
				RD_ADD(1), "RAD1",
				0.0 ns,
				RD_CLK, "RCLK",
				0.0 ns,
				tsetup_RAD1_RCLK_noedge_posedge, tsetup_RAD1_RCLK_noedge_posedge, 
				thold_RAD1_RCLK_noedge_posedge, thold_RAD1_RCLK_noedge_posedge,
				REN_ipd = '1' ,
				'/',
				InstancePath & "/R_SS",
				TRUE,
				TRUE,
				WARNING );

	VitalSetupHoldCheck    (Tviol_RD_ADD_stp_hld_2,
				TimingData_RD_ADD_stp_hld_2,
				RD_ADD(2), "RAD2",
				0.0 ns,
				RD_CLK, "RCLK",
				0.0 ns,
				tsetup_RAD2_RCLK_noedge_posedge, tsetup_RAD2_RCLK_noedge_posedge, 
				thold_RAD2_RCLK_noedge_posedge, thold_RAD2_RCLK_noedge_posedge,
				REN_ipd = '1' ,
				'/',
				InstancePath & "/R_SS",
				TRUE,
				TRUE,
				WARNING );

	VitalSetupHoldCheck    (Tviol_RD_ADD_stp_hld_3,
				TimingData_RD_ADD_stp_hld_3,
				RD_ADD(3), "RAD3",
				0.0 ns,
				RD_CLK, "RCLK",
				0.0 ns,
				tsetup_RAD3_RCLK_noedge_posedge, tsetup_RAD3_RCLK_noedge_posedge, 
				thold_RAD3_RCLK_noedge_posedge, thold_RAD3_RCLK_noedge_posedge,
				REN_ipd = '1' ,
				'/',
				InstancePath & "/R_SS",
				TRUE,
				TRUE,
				WARNING );

	VitalSetupHoldCheck    (Tviol_RD_ADD_stp_hld_4,
				TimingData_RD_ADD_stp_hld_4,
				RD_ADD(4), "RAD4",
				0.0 ns,
				RD_CLK, "RCLK",
				0.0 ns,
				tsetup_RAD4_RCLK_noedge_posedge, tsetup_RAD4_RCLK_noedge_posedge, 
				thold_RAD4_RCLK_noedge_posedge, thold_RAD4_RCLK_noedge_posedge,
				REN_ipd = '1' ,
				'/',
				InstancePath & "/R_SS",
				TRUE,
				TRUE,
				WARNING );

	VitalSetupHoldCheck    (Tviol_REN_hld,
				TimingData_REN_hld,
				REN_ipd, "REN",
				0.0 ns,
				RD_CLK, "RCLK",
				0.0 ns,
				tsetup_REN_RCLK_noedge_posedge, tsetup_REN_RCLK_noedge_posedge,
				thold_REN_RCLK_noedge_posedge, thold_REN_RCLK_noedge_posedge,
				True,
				'/',
				InstancePath & "/R_SS",
				TRUE,
				TRUE,
				WARNING );

    END IF; -- Timing Check Section

    -------------------------------------------------------------------
    -- Functionality Section
    -------------------------------------------------------------------

if (first) then
          while( not(endfile(STF)) ) loop
                readline(STF,readdata) ;
                read(readdata,tmp_data) ;
                memory_array(T) := tmp_data;
                T := T + 1;
              end loop;
end if;


-- READ ADDRESS CYCLE VIOLATION EFFECT

    if( Tviol_RD_ADD_stp_hld_0 = 'X' or Tviol_RD_ADD_stp_hld_1 = 'X' or Tviol_RD_ADD_stp_hld_2 = 'X' or Tviol_RD_ADD_stp_hld_3 = 'X' or Tviol_RD_ADD_stp_hld_4 = 'X' or Pviol_RCLK = 'X' or Tviol_REN_hld = 'X' or (RD_CLK'EVENT and RD_CLK = '1' and vecX(RD_ADD))) then
	--output_delay <= 0 ns;
	data_out <= x_data;
    elsif

-- VALID MEMORY READ

    (RD_CLK'EVENT and RD_CLK = '1' and not( Tviol_RD_ADD_stp_hld_0 = 'X' or Tviol_RD_ADD_stp_hld_1 = 'X' or Tviol_RD_ADD_stp_hld_2 = 'X' or Tviol_RD_ADD_stp_hld_3 = 'X' or Tviol_RD_ADD_stp_hld_4 = 'X' or Pviol_RCLK = 'X' or Tviol_REN_hld = 'X' or vecX(RD_ADD)) ) then
	rd_address := vec2int(RD_ADD);
	--output_delay <= tpd_RCLK_RDATA_posedge(0);
	data_out <= memory_array(rd_address);
    end if;

    if RD_CLK'EVENT and RD_CLK /= RCLK_ipd and RD_CLK'LAST_VALUE = '1' then
	--output_delay <= 0 ns;
	data_out <= x_data;
    end if;


  END PROCESS;

    -------------------------------------------------------------------------------
    -- Temporary output signal should get assigned to the output signal.
    -------------------------------------------------------------------------------

    --RDATA <= data_out after output_delay;

   PROCESS(data_out, RCLK_ipd)

      VARIABLE GLITCH : VitalGlitchDataType;
      VARIABLE RDATA3_1 : std_logic := 'X';
      VARIABLE RDATA2_1 : std_logic := 'X';
      VARIABLE RDATA1_1 : std_logic := 'X';
      VARIABLE RDATA0_1 : std_logic := 'X';
     
   BEGIN
       RDATA3_1 := VitalBUF(data_out(3));
       RDATA2_1 := VitalBUF(data_out(2));
       RDATA1_1 := VitalBUF(data_out(1));
       RDATA0_1 := VitalBUF(data_out(0));

     VitalPathDelay01 ( RDATA3, GLITCH, "RDATA3", RDATA3_1,
        Paths => (
        0 => ( RCLK_ipd'LAST_EVENT, tpd_RCLK_RDATA3, TRUE )),
        DefaultDelay=>VitalZeroDelay01,
        Mode=>VitalInertial,
        XON=>TRUE,
        MsgOn=>TRUE,
        MsgSeverity=>WARNING );

     VitalPathDelay01 ( RDATA2, GLITCH, "RDATA2", RDATA2_1,
        Paths => (
        0 => ( RCLK_ipd'LAST_EVENT, tpd_RCLK_RDATA2, TRUE )),
        DefaultDelay=>VitalZeroDelay01,
        Mode=>VitalInertial,
        XON=>TRUE,
        MsgOn=>TRUE,
        MsgSeverity=>WARNING );

     VitalPathDelay01 ( RDATA1, GLITCH, "RDATA1", RDATA1_1,
        Paths => (
        0 => ( RCLK_ipd'LAST_EVENT, tpd_RCLK_RDATA1, TRUE )),
        DefaultDelay=>VitalZeroDelay01,
        Mode=>VitalInertial,
        XON=>TRUE,
        MsgOn=>TRUE,
        MsgSeverity=>WARNING );

     VitalPathDelay01 ( RDATA0, GLITCH, "RDATA0", RDATA0_1,
        Paths => (
        0 => ( RCLK_ipd'LAST_EVENT, tpd_RCLK_RDATA0, TRUE )),
        DefaultDelay=>VitalZeroDelay01,
        Mode=>VitalInertial,
        XON=>TRUE,
        MsgOn=>TRUE,
        MsgSeverity=>WARNING );

END PROCESS;

END VITAL_VF;
configuration CFG_R_SS_VITAL of R_SS is
        for VITAL_VF
        end for;
end CFG_R_SS_VITAL;
-----------------------------------------------------------------------

----------------------------------------------------------------------- 
-- VITAL model for R_DAR 30.10 technology 
----------------------------------------------------------------------- 
 
LIBRARY IEEE; 
USE IEEE.std_logic_1164.ALL; 
USE IEEE.VITAL_timing.all; 
USE IEEE.std_logic_textio.all; 
USE IEEE.VITAL_primitives.all; 
LIBRARY std; 
USE std.textio.all; 
LIBRARY VF1; 
USE VF1.ALL; 
USE VF1.RAMPACK.ALL; 
 
----------------------------------------------------------------------- 
-- ENTITY declaration 
----------------------------------------------------------------------- 
 
ENTITY R_DAR IS 
  GENERIC ( 
	tipd_REN		: VitalDelayType01			:= (0.0 ns, 0.0 ns); 
	tipd_OE			: VitalDelayType01			:= (0.0 ns, 0.0 ns); 
	tipd_ADRCLK		: VitalDelayType01			:= (0.0 ns, 0.0 ns); 
	tipd_RAD10		: VitalDelayType01			:= (0.0 ns, 0.0 ns); 
	tipd_RAD11		: VitalDelayType01			:= (0.0 ns, 0.0 ns); 
	tipd_RAD12		: VitalDelayType01			:= (0.0 ns, 0.0 ns); 
	tipd_RAD13		: VitalDelayType01			:= (0.0 ns, 0.0 ns); 
	tipd_RAD14		: VitalDelayType01			:= (0.0 ns, 0.0 ns); 
	tipd_RAD20		: VitalDelayType01			:= (0.0 ns, 0.0 ns); 
	tipd_RAD21		: VitalDelayType01			:= (0.0 ns, 0.0 ns); 
	tipd_RAD22		: VitalDelayType01			:= (0.0 ns, 0.0 ns); 
	tipd_RAD23		: VitalDelayType01			:= (0.0 ns, 0.0 ns); 
	tipd_RAD24		: VitalDelayType01			:= (0.0 ns, 0.0 ns); 
 
tpd_ADRCLK_RDATA20         :VitalDelayType01 := (2.0 ns,2.0 ns);
tpd_ADRCLK_RDATA21         :VitalDelayType01 := (2.0 ns,2.0 ns);
tpd_ADRCLK_RDATA22         :VitalDelayType01 := (2.0 ns,2.0 ns);
tpd_ADRCLK_RDATA23         :VitalDelayType01 := (2.0 ns,2.0 ns);
tpd_OE_RDATA20         :VitalDelayType01 := (2.0 ns,2.0 ns);
tpd_OE_RDATA21         :VitalDelayType01 := (2.0 ns,2.0 ns);
tpd_OE_RDATA22         :VitalDelayType01 := (2.0 ns,2.0 ns);
tpd_OE_RDATA23         :VitalDelayType01 := (2.0 ns,2.0 ns);
tpd_ADRCLK_RDATA10         :VitalDelayType01 := (2.0 ns,2.0 ns);
tpd_ADRCLK_RDATA11         :VitalDelayType01 := (2.0 ns,2.0 ns);
tpd_ADRCLK_RDATA12         :VitalDelayType01 := (2.0 ns,2.0 ns);
tpd_ADRCLK_RDATA13         :VitalDelayType01 := (2.0 ns,2.0 ns);
tpw_ADRCLK_posedge        :VitalDelayType := 1.0 ns;

 
	tsetup_RAD10_ADRCLK_noedge_posedge		: VitalDelayType := 1 ns; 
	tsetup_RAD11_ADRCLK_noedge_posedge		: VitalDelayType := 1 ns; 
	tsetup_RAD12_ADRCLK_noedge_posedge		: VitalDelayType := 1 ns; 
	tsetup_RAD13_ADRCLK_noedge_posedge		: VitalDelayType := 1 ns; 
	tsetup_RAD14_ADRCLK_noedge_posedge		: VitalDelayType := 1 ns; 
	thold_RAD10_ADRCLK_noedge_posedge		: VitalDelayType := 1 ns; 
	thold_RAD11_ADRCLK_noedge_posedge		: VitalDelayType := 1 ns; 
	thold_RAD12_ADRCLK_noedge_posedge		: VitalDelayType := 1 ns; 
	thold_RAD13_ADRCLK_noedge_posedge		: VitalDelayType := 1 ns; 
	thold_RAD14_ADRCLK_noedge_posedge		: VitalDelayType := 1 ns; 

	tsetup_RAD20_ADRCLK_noedge_posedge		: VitalDelayType := 1 ns; 
	tsetup_RAD21_ADRCLK_noedge_posedge		: VitalDelayType := 1 ns; 
	tsetup_RAD22_ADRCLK_noedge_posedge		: VitalDelayType := 1 ns; 
	tsetup_RAD23_ADRCLK_noedge_posedge		: VitalDelayType := 1 ns; 
	tsetup_RAD24_ADRCLK_noedge_posedge		: VitalDelayType := 1 ns; 
	thold_RAD20_ADRCLK_noedge_posedge		: VitalDelayType := 1 ns; 
	thold_RAD21_ADRCLK_noedge_posedge		: VitalDelayType := 1 ns; 
	thold_RAD22_ADRCLK_noedge_posedge		: VitalDelayType := 1 ns; 
	thold_RAD23_ADRCLK_noedge_posedge		: VitalDelayType := 1 ns; 
	thold_RAD24_ADRCLK_noedge_posedge		: VitalDelayType := 1 ns; 

 
	TimingChecksOn : BOOLEAN := TRUE; 
	InstancePath : STRING := "*" 
            ); 
  PORT	( 
	REN		: IN	std_logic ; 
	OE		: IN	std_logic ; 
	ADRCLK		: IN	std_logic ; 
	RDATA20	        : OUT	std_logic := 'X'; 
	RDATA21	        : OUT	std_logic := 'X'; 
	RDATA22	        : OUT	std_logic := 'X'; 
	RDATA23	        : OUT	std_logic := 'X'; 
	RDATA10		: OUT	std_logic := 'X'; 
	RDATA11		: OUT	std_logic := 'X'; 
	RDATA12		: OUT	std_logic := 'X'; 
	RDATA13		: OUT	std_logic := 'X'; 
	RAD10		: IN	std_logic; 
	RAD11		: IN	std_logic; 
	RAD12		: IN	std_logic; 
	RAD13		: IN	std_logic; 
	RAD14		: IN	std_logic; 
	RAD20		: IN	std_logic; 
	RAD21		: IN	std_logic; 
	RAD22		: IN	std_logic; 
	RAD23		: IN	std_logic; 
	RAD24		: IN	std_logic 
	); 
 
 
   ATTRIBUTE VITAL_LEVEL0 OF R_DAR : ENTITY IS TRUE; 
 
END R_DAR; 
 
----------------------------------------------------------------------- 
-- ARCHITECTURE declaration 
----------------------------------------------------------------------- 
ARCHITECTURE VITAL_VF OF R_DAR IS 
 
    ATTRIBUTE VITAL_LEVEL1 OF VITAL_VF : ARCHITECTURE IS FALSE; 
 
	file STF : text is in "rom_data"; 
	SIGNAL REN_ipd		: std_logic := '0'; 
	SIGNAL OE_ipd	: std_logic := '0'; 
	SIGNAL ADRCLK_ipd	: std_logic := '0'; 
	SIGNAL RAD10_ipd		: std_logic; 
	SIGNAL RAD11_ipd		: std_logic; 
	SIGNAL RAD12_ipd		: std_logic; 
	SIGNAL RAD13_ipd		: std_logic; 
	SIGNAL RAD14_ipd		: std_logic; 
	SIGNAL RD_ADD1		: std_logic_vector(4 DOWNTO 0); 
	SIGNAL RD_ADD2		: std_logic_vector(4 DOWNTO 0); 
	SIGNAL RAD20_ipd		: std_logic; 
	SIGNAL RAD21_ipd		: std_logic; 
	SIGNAL RAD22_ipd		: std_logic; 
	SIGNAL RAD23_ipd		: std_logic; 
	SIGNAL RAD24_ipd		: std_logic; 
	SIGNAL data_out		: std_logic_vector(3 DOWNTO 0) := x_data; 
	SIGNAL data_out_w	: std_logic_vector(3 DOWNTO 0) := x_data; 
	SIGNAL output_delay	: time		:= 0 ns; 
	SIGNAL output_delay_w	: time		:= 0 ns; 
	SIGNAL memory_array	: memory_array_typ; 
 
BEGIN 
    
  --------------------------------------------------------------------- 
  -- INPUT PATH DELAYs 
  --------------------------------------------------------------------- 
  WIREDELAY : BLOCK 
  BEGIN 
	VitalWireDelay (REN_ipd,		REN,		tipd_REN); 
	VitalWireDelay (OE_ipd,		OE,		tipd_OE); 
	VitalWireDelay (ADRCLK_ipd,		ADRCLK,		tipd_ADRCLK); 
        VitalWireDelay (RAD10_ipd,              RAD10,          tipd_RAD10);
        VitalWireDelay (RAD11_ipd,              RAD11,          tipd_RAD11);
        VitalWireDelay (RAD12_ipd,              RAD12,          tipd_RAD12);
        VitalWireDelay (RAD13_ipd,              RAD13,          tipd_RAD13);
        VitalWireDelay (RAD14_ipd,              RAD14,          tipd_RAD14);
        VitalWireDelay (RAD20_ipd,              RAD20,          tipd_RAD20);
        VitalWireDelay (RAD21_ipd,              RAD21,          tipd_RAD21);
        VitalWireDelay (RAD22_ipd,              RAD22,          tipd_RAD22);
        VitalWireDelay (RAD23_ipd,              RAD23,          tipd_RAD23);
        VitalWireDelay (RAD24_ipd,              RAD24,          tipd_RAD24);

  END BLOCK; 
 
  --------------------------------------------------------------------- 
  -- Behavior Section 
  --------------------------------------------------------------------- 
 
  --------------------------------------------------------------------- 
  -- Wrapper Section 
  --------------------------------------------------------------------- 
 
   wrapper_latch_add : process(ADRCLK_ipd) 
 
   begin 
    if (ADRCLK_ipd = '1' ) then 
	RD_ADD1(4) <= RAD14_ipd; 
	RD_ADD1(3) <= RAD13_ipd; 
	RD_ADD1(2) <= RAD12_ipd; 
	RD_ADD1(1) <= RAD11_ipd; 
	RD_ADD1(0) <= RAD10_ipd; 
	RD_ADD2(4) <= RAD24_ipd; 
	RD_ADD2(3) <= RAD23_ipd; 
	RD_ADD2(2) <= RAD22_ipd; 
	RD_ADD2(1) <= RAD21_ipd; 
	RD_ADD2(0) <= RAD20_ipd; 
    end if; 
 
   end process; 
 
 
  VITALBehavior : PROCESS ( REN_ipd, OE_ipd, RD_ADD2, RD_ADD1, ADRCLK_ipd, RAD14_ipd, RAD13_ipd, RAD12_ipd, RAD11_ipd, RAD10_ipd, RAD24_ipd, RAD23_ipd, RAD22_ipd, RAD21_ipd, RAD20_ipd ) 
 
 
   -- Temporary variables 
   VARIABLE tmp_data : std_logic_vector (3 downto 0); 
   VARIABLE readdata : LINE; 
   VARIABLE first : boolean := TRUE; 
   VARIABLE rd_address 		: integer := 0; 
   VARIABLE rd_address_w 	: integer := 0; 
   VARIABLE T 	: integer := 0; 
   VARIABLE rd_viol_flag 	: X01 := '0'; 
   VARIABLE rd_viol_flag_w 	: X01 := '0'; 
 
   -- Timing Check results 
   VARIABLE Pviol_ADRCLK		: std_logic := '0'; 
   VARIABLE PeriodData_ADRCLK		: VitalPeriodDataType := VitalPeriodDataInit; 
   VARIABLE Tviol_RAD1_stp_hld_0		: std_logic := '0'; 
   VARIABLE TimingData_RAD1_stp_hld_0	: VitalTimingDataType := VitalTimingDataInit; 
   VARIABLE Tviol_RAD1_stp_hld_1		: std_logic := '0'; 
   VARIABLE TimingData_RAD1_stp_hld_1	: VitalTimingDataType := VitalTimingDataInit; 
   VARIABLE Tviol_RAD1_stp_hld_2		: std_logic := '0'; 
   VARIABLE TimingData_RAD1_stp_hld_2	: VitalTimingDataType := VitalTimingDataInit; 
   VARIABLE Tviol_RAD1_stp_hld_3		: std_logic := '0'; 
   VARIABLE TimingData_RAD1_stp_hld_3	: VitalTimingDataType := VitalTimingDataInit; 
   VARIABLE Tviol_RAD1_stp_hld_4		: std_logic := '0'; 
   VARIABLE TimingData_RAD1_stp_hld_4	: VitalTimingDataType := VitalTimingDataInit; 
   VARIABLE Tviol_RAD2_stp_hld_0		: std_logic := '0'; 
   VARIABLE TimingData_RAD2_stp_hld_0	: VitalTimingDataType := VitalTimingDataInit; 
   VARIABLE Tviol_RAD2_stp_hld_1		: std_logic := '0'; 
   VARIABLE TimingData_RAD2_stp_hld_1	: VitalTimingDataType := VitalTimingDataInit; 
   VARIABLE Tviol_RAD2_stp_hld_2		: std_logic := '0'; 
   VARIABLE TimingData_RAD2_stp_hld_2	: VitalTimingDataType := VitalTimingDataInit; 
   VARIABLE Tviol_RAD2_stp_hld_3		: std_logic := '0'; 
   VARIABLE TimingData_RAD2_stp_hld_3	: VitalTimingDataType := VitalTimingDataInit; 
   VARIABLE Tviol_RAD2_stp_hld_4		: std_logic := '0'; 
   VARIABLE TimingData_RAD2_stp_hld_4	: VitalTimingDataType := VitalTimingDataInit; 
 
 
 
 BEGIN 
    ------------------------------------------------------------------- 
    -- Timing Check Section 
    ------------------------------------------------------------------- 
    IF (TimingChecksOn) THEN 
 
	VitalPeriodPulseCheck  (Pviol_ADRCLK, 
				PeriodData_ADRCLK, 
				ADRCLK_ipd, "ADRCLK", 
				0.0 ns, 
				0.0 ns, 
				tpw_ADRCLK_posedge, 
				0.0 ns, 
				True ,
				InstancePath & "/R_DAR", 
				TRUE, 
				TRUE, 
				WARNING ); 
 
 
	VitalSetupHoldCheck    (Tviol_RAD1_stp_hld_0, 
				TimingData_RAD1_stp_hld_0, 
				RAD10_ipd, "RAD10", 
				0.0 ns, 
				ADRCLK_ipd, "ADRCLK", 
				0.0 ns, 
				tsetup_RAD10_ADRCLK_noedge_posedge,tsetup_RAD10_ADRCLK_noedge_posedge,
				thold_RAD10_ADRCLK_noedge_posedge,thold_RAD10_ADRCLK_noedge_posedge,
				REN_ipd = '1', 
				'/', 
				InstancePath & "/R_DAR", 
				TRUE, 
				TRUE, 
				WARNING ); 
 
	VitalSetupHoldCheck    (Tviol_RAD1_stp_hld_1, 
				TimingData_RAD1_stp_hld_1, 
				RAD11_ipd, "RAD11", 
				0.0 ns, 
				ADRCLK_ipd, "ADRCLK", 
				0.0 ns, 
				tsetup_RAD11_ADRCLK_noedge_posedge,tsetup_RAD11_ADRCLK_noedge_posedge,
				thold_RAD11_ADRCLK_noedge_posedge,thold_RAD11_ADRCLK_noedge_posedge,
				REN_ipd = '1', 
				'/', 
				InstancePath & "/R_DAR", 
				TRUE, 
				TRUE, 
				WARNING ); 
 
	VitalSetupHoldCheck    (Tviol_RAD1_stp_hld_2, 
				TimingData_RAD1_stp_hld_2, 
				RAD12_ipd, "RAD12", 
				0.0 ns, 
				ADRCLK_ipd, "ADRCLK", 
				0.0 ns, 
				tsetup_RAD12_ADRCLK_noedge_posedge,tsetup_RAD12_ADRCLK_noedge_posedge,
				thold_RAD12_ADRCLK_noedge_posedge,thold_RAD12_ADRCLK_noedge_posedge,
				REN_ipd = '1', 
				'/', 
				InstancePath & "/R_DAR", 
				TRUE, 
				TRUE, 
				WARNING ); 

	VitalSetupHoldCheck    (Tviol_RAD1_stp_hld_3, 
				TimingData_RAD1_stp_hld_3, 
				RAD13_ipd, "RAD13", 
				0.0 ns, 
				ADRCLK_ipd, "ADRCLK", 
				0.0 ns, 
				tsetup_RAD13_ADRCLK_noedge_posedge,tsetup_RAD13_ADRCLK_noedge_posedge,
				thold_RAD13_ADRCLK_noedge_posedge,thold_RAD13_ADRCLK_noedge_posedge,
				REN_ipd = '1', 
				'/', 
				InstancePath & "/R_DAR", 
				TRUE, 
				TRUE, 
				WARNING ); 

	VitalSetupHoldCheck    (Tviol_RAD1_stp_hld_4, 
				TimingData_RAD1_stp_hld_4, 
				RAD14_ipd, "RAD14", 
				0.0 ns, 
				ADRCLK_ipd, "ADRCLK", 
				0.0 ns, 
				tsetup_RAD14_ADRCLK_noedge_posedge,tsetup_RAD14_ADRCLK_noedge_posedge,
				thold_RAD14_ADRCLK_noedge_posedge,thold_RAD14_ADRCLK_noedge_posedge,
				REN_ipd = '1', 
				'/', 
				InstancePath & "/R_DAR", 
				TRUE, 
				TRUE, 
				WARNING ); 

	VitalSetupHoldCheck    (Tviol_RAD2_stp_hld_0, 
				TimingData_RAD2_stp_hld_0, 
				RAD20_ipd, "RAD20", 
				0.0 ns, 
				ADRCLK_ipd, "ADRCLK", 
				0.0 ns, 
				tsetup_RAD20_ADRCLK_noedge_posedge,tsetup_RAD20_ADRCLK_noedge_posedge,
				thold_RAD20_ADRCLK_noedge_posedge,thold_RAD20_ADRCLK_noedge_posedge,
				REN_ipd = '1', 
				'/', 
				InstancePath & "/R_DAR", 
				TRUE, 
				TRUE, 
				WARNING ); 
 
	VitalSetupHoldCheck    (Tviol_RAD2_stp_hld_1, 
				TimingData_RAD2_stp_hld_1, 
				RAD21_ipd, "RAD21", 
				0.0 ns, 
				ADRCLK_ipd, "ADRCLK", 
				0.0 ns, 
				tsetup_RAD21_ADRCLK_noedge_posedge,tsetup_RAD21_ADRCLK_noedge_posedge,
				thold_RAD21_ADRCLK_noedge_posedge,thold_RAD21_ADRCLK_noedge_posedge,
				REN_ipd = '1', 
				'/', 
				InstancePath & "/R_DAR", 
				TRUE, 
				TRUE, 
				WARNING ); 
 
	VitalSetupHoldCheck    (Tviol_RAD2_stp_hld_2, 
				TimingData_RAD2_stp_hld_2, 
				RAD22_ipd, "RAD22", 
				0.0 ns, 
				ADRCLK_ipd, "ADRCLK", 
				0.0 ns, 
				tsetup_RAD22_ADRCLK_noedge_posedge,tsetup_RAD22_ADRCLK_noedge_posedge,
				thold_RAD22_ADRCLK_noedge_posedge,thold_RAD22_ADRCLK_noedge_posedge,
				REN_ipd = '1', 
				'/', 
				InstancePath & "/R_DAR", 
				TRUE, 
				TRUE, 
				WARNING ); 

	VitalSetupHoldCheck    (Tviol_RAD2_stp_hld_3, 
				TimingData_RAD2_stp_hld_3, 
				RAD23_ipd, "RAD23", 
				0.0 ns, 
				ADRCLK_ipd, "ADRCLK", 
				0.0 ns, 
				tsetup_RAD23_ADRCLK_noedge_posedge,tsetup_RAD23_ADRCLK_noedge_posedge,
				thold_RAD23_ADRCLK_noedge_posedge,thold_RAD23_ADRCLK_noedge_posedge,
				REN_ipd = '1', 
				'/', 
				InstancePath & "/R_DAR", 
				TRUE, 
				TRUE, 
				WARNING ); 

	VitalSetupHoldCheck    (Tviol_RAD2_stp_hld_4, 
				TimingData_RAD2_stp_hld_4, 
				RAD24_ipd, "RAD24", 
				0.0 ns, 
				ADRCLK_ipd, "ADRCLK", 
				0.0 ns, 
				tsetup_RAD24_ADRCLK_noedge_posedge,tsetup_RAD24_ADRCLK_noedge_posedge,
				thold_RAD24_ADRCLK_noedge_posedge,thold_RAD24_ADRCLK_noedge_posedge,
				REN_ipd = '1', 
				'/', 
				InstancePath & "/R_DAR", 
				TRUE, 
				TRUE, 
                                WARNING );


    END IF; -- Timing Check Section 
 
rd_viol_flag := (Tviol_RAD1_stp_hld_0 or Tviol_RAD1_stp_hld_1 or Tviol_RAD1_stp_hld_2 or Tviol_RAD1_stp_hld_3 or Tviol_RAD1_stp_hld_4 or Pviol_ADRCLK ); 

rd_viol_flag_w := (Tviol_RAD2_stp_hld_0 or Tviol_RAD2_stp_hld_1 or Tviol_RAD2_stp_hld_2 or Tviol_RAD2_stp_hld_3 or Tviol_RAD2_stp_hld_4 or Pviol_ADRCLK ); 
 
 
 
 
    ------------------------------------------------------------------- 
    -- Functionality Section 
    ------------------------------------------------------------------- 
 
 
if (first) then 
          while( not(endfile(STF)) ) loop 
                readline(STF,readdata) ; 
                read(readdata,tmp_data) ; 
 
  --for T in 0 to 31 loop 
   -- READLINE (STF,readdata); 
    --Read (readdata,tmp_data); 
    memory_array(T) <= tmp_data; 
   T := T + 1; 
  end loop; 
   first := FALSE;
end if; 
 
 
 
-- READ CYCLE VIOLATION EFFECT 
 
    if( rd_viol_flag = 'X'  or (RD_ADD1'EVENT  and REN_ipd = '1' and vecX(RD_ADD1))) then 
	--output_delay <= 0 ns; 
	data_out <= x_data; 
    elsif 
 
-- VALID MEMORY READ 
 
 
     (RD_ADD1'EVENT and REN_ipd = '1' and not(rd_viol_flag = 'X') and not (vecX(RD_ADD1))) then 
	rd_address := vec2int(RD_ADD1); 
	data_out <= memory_array(rd_address); 
    end if; 
 
 
    if( rd_viol_flag_w = 'X' or (RD_ADD2'EVENT and REN_ipd = '1' and OE_ipd = '1' and vecX(RD_ADD2))) then 
	--output_delay_w <= 0 ns; 
	data_out_w <= x_data; 
    elsif 
 
-- VALID MEMORY READ 
 
     (RD_ADD2'EVENT and REN_ipd = '1' and OE_ipd = '1'  and not(rd_viol_flag_w = 'X') and not (vecX(RD_ADD2))) then 
	rd_address_w := vec2int(RD_ADD2); 
	data_out_w <= memory_array(rd_address_w); 
    end if; 
 
 
  END PROCESS; 
 
    ------------------------------------------------------------------------------- 
    -- Temporary output signal should get assigned to the output signal. 
    ------------------------------------------------------------------------------- 
 
   -- RDATA1 <= TRANSPORT data_out after output_delay; 
 
 
   PROCESS(data_out, data_out_w, ADRCLK_ipd, OE_ipd)

      VARIABLE GLITCH1 : VitalGlitchDataType;
      VARIABLE GLITCH2 : VitalGlitchDataType;
      VARIABLE RDATA13_1 : std_logic := 'X';
      VARIABLE RDATA12_1 : std_logic := 'X';
      VARIABLE RDATA11_1 : std_logic := 'X';
      VARIABLE RDATA10_1 : std_logic := 'X';
      VARIABLE RDATA23_1 : std_logic := 'X';
      VARIABLE RDATA22_1 : std_logic := 'X';
      VARIABLE RDATA21_1 : std_logic := 'X';
      VARIABLE RDATA20_1 : std_logic := 'X';

   BEGIN
       RDATA23_1 := VitalBUF(data_out_w(3));
       RDATA22_1 := VitalBUF(data_out_w(2));
       RDATA21_1 := VitalBUF(data_out_w(1));
       RDATA20_1 := VitalBUF(data_out_w(0));
       RDATA13_1 := VitalBUF(data_out(3));
       RDATA12_1 := VitalBUF(data_out(2));
       RDATA11_1 := VitalBUF(data_out(1));
       RDATA10_1 := VitalBUF(data_out(0));

     VitalPathDelay01 ( RDATA13, GLITCH1, "RDATA13", RDATA13_1,
        Paths => (
        0 => ( ADRCLK_ipd'LAST_EVENT, tpd_ADRCLK_RDATA13, TRUE )),
        DefaultDelay=>VitalZeroDelay01,
        Mode=>VitalInertial,
        XON=>TRUE,
        MsgOn=>TRUE,
        MsgSeverity=>WARNING );

     VitalPathDelay01 ( RDATA12, GLITCH1, "RDATA12", RDATA12_1,
        Paths => (
        0 => ( ADRCLK_ipd'LAST_EVENT, tpd_ADRCLK_RDATA12, TRUE )),
        DefaultDelay=>VitalZeroDelay01,
        Mode=>VitalInertial,
        XON=>TRUE,
        MsgOn=>TRUE,
        MsgSeverity=>WARNING );

     VitalPathDelay01 ( RDATA11, GLITCH1, "RDATA11", RDATA11_1,
        Paths => (
        0 => ( ADRCLK_ipd'LAST_EVENT, tpd_ADRCLK_RDATA11, TRUE )),
        DefaultDelay=>VitalZeroDelay01,
        Mode=>VitalInertial,
        XON=>TRUE,
        MsgOn=>TRUE,
        MsgSeverity=>WARNING );

     VitalPathDelay01 ( RDATA10, GLITCH1, "RDATA10", RDATA10_1,
        Paths => (
        0 => ( ADRCLK_ipd'LAST_EVENT, tpd_ADRCLK_RDATA10, TRUE )),
        DefaultDelay=>VitalZeroDelay01,
        Mode=>VitalInertial,
        XON=>TRUE,
        MsgOn=>TRUE,
        MsgSeverity=>WARNING );

     VitalPathDelay01 ( RDATA23, GLITCH2, "RDATA23", RDATA23_1,
        Paths => (
        0 => ( ADRCLK_ipd'LAST_EVENT, tpd_ADRCLK_RDATA23, TRUE ),
        1 => ( OE_ipd'LAST_EVENT, tpd_OE_RDATA23, TRUE )),
        DefaultDelay=>VitalZeroDelay01,
        Mode=>VitalInertial,
        XON=>TRUE,
        MsgOn=>TRUE,
        MsgSeverity=>WARNING );

     VitalPathDelay01 ( RDATA22, GLITCH2, "RDATA22", RDATA22_1,
        Paths => (
        0 => ( ADRCLK_ipd'LAST_EVENT, tpd_ADRCLK_RDATA22, TRUE ),
        1 => ( OE_ipd'LAST_EVENT, tpd_OE_RDATA22, TRUE )),
        DefaultDelay=>VitalZeroDelay01,
        Mode=>VitalInertial,
        XON=>TRUE,
        MsgOn=>TRUE,
        MsgSeverity=>WARNING );

     VitalPathDelay01 ( RDATA21, GLITCH2, "RDATA21", RDATA21_1,
        Paths => (
        0 => ( ADRCLK_ipd'LAST_EVENT, tpd_ADRCLK_RDATA21, TRUE ),
        1 => ( OE_ipd'LAST_EVENT, tpd_OE_RDATA21, TRUE )),
        DefaultDelay=>VitalZeroDelay01,
        Mode=>VitalInertial,
        XON=>TRUE,
        MsgOn=>TRUE,
        MsgSeverity=>WARNING );

     VitalPathDelay01 ( RDATA20, GLITCH2, "RDATA20", RDATA20_1,
        Paths => (
        0 => ( ADRCLK_ipd'LAST_EVENT, tpd_ADRCLK_RDATA20, TRUE ),
        1 => ( OE_ipd'LAST_EVENT, tpd_OE_RDATA20, TRUE )),
        DefaultDelay=>VitalZeroDelay01,
        Mode=>VitalInertial,
        XON=>TRUE,
        MsgOn=>TRUE,
        MsgSeverity=>WARNING );

END PROCESS;
 
END VITAL_VF; 
configuration CFG_R_DAR_VITAL of R_DAR is
        for VITAL_VF
        end for;
end CFG_R_DAR_VITAL;
 
-----------------------------------------------------------------------
-- VITAL model for R_SAR 30.10 technology 
----------------------------------------------------------------------- 
 
LIBRARY IEEE; 
USE IEEE.std_logic_1164.ALL; 
USE IEEE.VITAL_timing.all; 
USE IEEE.VITAL_primitives.all; 
USE IEEE.std_logic_textio.all; 
LIBRARY std; 
USE std.textio.all; 
LIBRARY VF1; 
USE VF1.ALL; 
USE VF1.RAMPACK.ALL; 
 
----------------------------------------------------------------------- 
-- ENTITY declaration 
----------------------------------------------------------------------- 
 
ENTITY R_SAR IS 
  GENERIC ( 
	tipd_REN		: VitalDelayType01			:= (0.0 ns, 0.0 ns); 
	tipd_ADRCLK		: VitalDelayType01			:= (0.0 ns, 0.0 ns); 
	tipd_RAD0		: VitalDelayType01	:= (0.0 ns, 0.0 ns); 
	tipd_RAD1		: VitalDelayType01	:= (0.0 ns, 0.0 ns); 
	tipd_RAD2		: VitalDelayType01	:= (0.0 ns, 0.0 ns); 
	tipd_RAD3		: VitalDelayType01	:= (0.0 ns, 0.0 ns); 
	tipd_RAD4		: VitalDelayType01	:= (0.0 ns, 0.0 ns); 
 
        tpd_ADRCLK_RDATA0                 : VitalDelayType01 := (2 ns,2 ns);
        tpd_ADRCLK_RDATA1                 : VitalDelayType01 := (2 ns,2 ns);
        tpd_ADRCLK_RDATA2                 : VitalDelayType01 := (2 ns,2 ns);
        tpd_ADRCLK_RDATA3                 : VitalDelayType01 := (2 ns,2 ns);

        tpd_REN_RDATA0                 : VitalDelayType01 := (2 ns,2 ns);
        tpd_REN_RDATA1                 : VitalDelayType01 := (2 ns,2 ns);
        tpd_REN_RDATA2                 : VitalDelayType01 := (2 ns,2 ns);
        tpd_REN_RDATA3                 : VitalDelayType01 := (2 ns,2 ns);



	tsetup_RAD0_ADRCLK_noedge_posedge	: VitalDelayType := 1 ns; 
	tsetup_RAD1_ADRCLK_noedge_posedge	: VitalDelayType := 1 ns; 
	tsetup_RAD2_ADRCLK_noedge_posedge	: VitalDelayType := 1 ns; 
	tsetup_RAD3_ADRCLK_noedge_posedge	: VitalDelayType := 1 ns; 
	tsetup_RAD4_ADRCLK_noedge_posedge	: VitalDelayType := 1 ns; 


	thold_RAD0_ADRCLK_noedge_posedge	: VitalDelayType := 1 ns; 
	thold_RAD1_ADRCLK_noedge_posedge	: VitalDelayType := 1 ns; 
	thold_RAD2_ADRCLK_noedge_posedge	: VitalDelayType := 1 ns; 
	thold_RAD3_ADRCLK_noedge_posedge	: VitalDelayType := 1 ns; 
	thold_RAD4_ADRCLK_noedge_posedge	: VitalDelayType := 1 ns; 

        tpw_ADRCLK_posedge                              : VitalDelayType := 1 ns;


	TimingChecksOn : BOOLEAN := TRUE; 
	InstancePath : STRING := "*" 
            ); 
  PORT	( 
	REN		: IN	std_logic ; 
	ADRCLK		: IN	std_logic ; 
	RDATA0		: OUT	std_logic := 'X'; 
	RDATA1		: OUT	std_logic := 'X'; 
	RDATA2		: OUT	std_logic := 'X'; 
	RDATA3		: OUT	std_logic := 'X'; 
	RAD0		: IN	std_logic;
	RAD1		: IN	std_logic;
	RAD2		: IN	std_logic;
	RAD3		: IN	std_logic;
	RAD4		: IN	std_logic 
	); 
 
 
   ATTRIBUTE VITAL_LEVEL0 OF R_SAR : ENTITY IS TRUE; 
 
END R_SAR; 
 
----------------------------------------------------------------------- 
-- ARCHITECTURE declaration 
----------------------------------------------------------------------- 
ARCHITECTURE VITAL_VF OF R_SAR IS 
 
    ATTRIBUTE VITAL_LEVEL1 OF VITAL_VF : ARCHITECTURE IS FALSE; 
 
	file STF : text is in "rom_data"; 
	SIGNAL REN_ipd		: std_logic := 'X'; 
	SIGNAL ADRCLK_ipd		: std_logic := '0'; 
	SIGNAL RAD0_ipd		: std_logic; 
	SIGNAL RAD1_ipd		: std_logic; 
	SIGNAL RAD2_ipd		: std_logic; 
	SIGNAL RAD3_ipd		: std_logic; 
	SIGNAL RAD4_ipd		: std_logic; 
	SIGNAL RD_ADD		: std_logic_vector(4 DOWNTO 0); 
	SIGNAL data_out		: std_logic_vector(3 DOWNTO 0) := x_data; 
	SIGNAL output_delay	: time		:= 0 ns; 
	SIGNAL memory_array	: memory_array_typ; 
 
BEGIN 
    
  --------------------------------------------------------------------- 
  -- INPUT PATH DELAYs 
  --------------------------------------------------------------------- 
  WIREDELAY : BLOCK 
  BEGIN 
	VitalWireDelay (REN_ipd,		REN,		tipd_REN); 
	VitalWireDelay (ADRCLK_ipd,		ADRCLK,		tipd_ADRCLK); 
	VitalWireDelay (RAD0_ipd,		RAD0,		tipd_RAD0); 
	VitalWireDelay (RAD1_ipd,		RAD1,		tipd_RAD1); 
	VitalWireDelay (RAD2_ipd,		RAD2,		tipd_RAD2); 
	VitalWireDelay (RAD3_ipd,		RAD3,		tipd_RAD3); 
	VitalWireDelay (RAD4_ipd,		RAD4,		tipd_RAD4); 
 
  END BLOCK; 
 
  --------------------------------------------------------------------- 
  -- Behavior Section 
  --------------------------------------------------------------------- 
 
  --------------------------------------------------------------------- 
  -- Wrapper Section 
  --------------------------------------------------------------------- 
 
   wrapper_latch_add : process(ADRCLK_ipd)--,RAD0_ipd,RAD1_ipd,RAD2_ipd,RAD3_ipd,RAD4_ipd) 
 
   begin 
    if (ADRCLK_ipd'EVENT and ADRCLK_ipd = '1' ) then 
	RD_ADD(0) <= RAD0_ipd; 
	RD_ADD(1) <= RAD1_ipd; 
	RD_ADD(2) <= RAD2_ipd; 
	RD_ADD(3) <= RAD3_ipd; 
	RD_ADD(4) <= RAD4_ipd; 
    end if; 
 
   end process; 
 
 
  VITALBehavior : PROCESS ( REN_ipd, ADRCLK_ipd, RD_ADD,  RAD0_ipd,  RAD1_ipd,  RAD2_ipd,  RAD3_ipd,  RAD4_ipd ) 
 
 
   -- Temporary variables 
   VARIABLE tmp_data : std_logic_vector (3 downto 0); 
   VARIABLE readdata : LINE; 
   VARIABLE first : boolean := TRUE; 
   VARIABLE rd_address 		: integer := 0; 
   VARIABLE T 		: integer := 0; 
   VARIABLE rd_viol_flag 	: X01 := '0'; 
 
   -- Timing Check results 
   VARIABLE Pviol_ADRCLK			: std_logic := '0'; 
   VARIABLE PeriodData_ADRCLK		: VitalPeriodDataType := VitalPeriodDataInit; 
   VARIABLE Tviol_RAD_stp_hld_0		: std_logic := '0'; 
   VARIABLE TimingData_RAD_stp_hld_0	: VitalTimingDataType := VitalTimingDataInit; 
   VARIABLE Tviol_RAD_stp_hld_1		: std_logic := '0'; 
   VARIABLE TimingData_RAD_stp_hld_1	: VitalTimingDataType := VitalTimingDataInit; 
   VARIABLE Tviol_RAD_stp_hld_2		: std_logic := '0'; 
   VARIABLE TimingData_RAD_stp_hld_2	: VitalTimingDataType := VitalTimingDataInit; 
   VARIABLE Tviol_RAD_stp_hld_3		: std_logic := '0'; 
   VARIABLE TimingData_RAD_stp_hld_3	: VitalTimingDataType := VitalTimingDataInit; 
   VARIABLE Tviol_RAD_stp_hld_4		: std_logic := '0'; 
   VARIABLE TimingData_RAD_stp_hld_4	: VitalTimingDataType := VitalTimingDataInit; 
 
 
 
 BEGIN 
    ------------------------------------------------------------------- 
    -- Timing Check Section 
    ------------------------------------------------------------------- 
    IF (TimingChecksOn) THEN 
 
	VitalPeriodPulseCheck  (Pviol_ADRCLK, 
				PeriodData_ADRCLK, 
				ADRCLK, "ADRCLK", 
				0.0 ns, 
				0.0 ns, 
				tpw_ADRCLK_posedge, 
				0.0 ns,
				True,
				InstancePath & "/R_SAR", 
				TRUE, 
				TRUE, 
				WARNING ); 
 
	VitalSetupHoldCheck    (Tviol_RAD_stp_hld_0, 
				TimingData_RAD_stp_hld_0, 
				RAD0_ipd, "RAD0", 
				0.0 ns, 
				ADRCLK_ipd, "ADRCLK", 
				0.0 ns, 
				tsetup_RAD0_ADRCLK_noedge_posedge, tsetup_RAD0_ADRCLK_noedge_posedge,
				thold_RAD0_ADRCLK_noedge_posedge, thold_RAD0_ADRCLK_noedge_posedge,
				REN_ipd = '1', 
				'/', 
				InstancePath & "/R_SAR", 
				TRUE, 
				TRUE, 
				WARNING ); 

	VitalSetupHoldCheck    (Tviol_RAD_stp_hld_1, 
				TimingData_RAD_stp_hld_1, 
				RAD1_ipd, "RAD1", 
				0.0 ns, 
				ADRCLK_ipd, "ADRCLK", 
				0.0 ns, 
				tsetup_RAD1_ADRCLK_noedge_posedge, tsetup_RAD1_ADRCLK_noedge_posedge,
				thold_RAD1_ADRCLK_noedge_posedge, thold_RAD1_ADRCLK_noedge_posedge,
				REN_ipd = '1', 
				'/', 
				InstancePath & "/R_SAR", 
				TRUE, 
				TRUE, 
				WARNING ); 

	VitalSetupHoldCheck    (Tviol_RAD_stp_hld_2, 
				TimingData_RAD_stp_hld_2, 
				RAD2_ipd, "RAD2", 
				0.0 ns, 
				ADRCLK_ipd, "ADRCLK", 
				0.0 ns, 
				tsetup_RAD2_ADRCLK_noedge_posedge, tsetup_RAD2_ADRCLK_noedge_posedge,
				thold_RAD2_ADRCLK_noedge_posedge, thold_RAD2_ADRCLK_noedge_posedge,
				REN_ipd = '1', 
				'/', 
				InstancePath & "/R_SAR", 
				TRUE, 
				TRUE, 
				WARNING ); 

	VitalSetupHoldCheck    (Tviol_RAD_stp_hld_3, 
				TimingData_RAD_stp_hld_3, 
				RAD3_ipd, "RAD3", 
				0.0 ns, 
				ADRCLK_ipd, "ADRCLK", 
				0.0 ns, 
				tsetup_RAD3_ADRCLK_noedge_posedge, tsetup_RAD3_ADRCLK_noedge_posedge,
				thold_RAD3_ADRCLK_noedge_posedge, thold_RAD3_ADRCLK_noedge_posedge,
				REN_ipd = '1', 
				'/', 
				InstancePath & "/R_SAR", 
				TRUE, 
				TRUE, 
				WARNING ); 

	VitalSetupHoldCheck    (Tviol_RAD_stp_hld_4, 
				TimingData_RAD_stp_hld_4, 
				RAD4_ipd, "RAD4", 
				0.0 ns, 
				ADRCLK_ipd, "ADRCLK", 
				0.0 ns, 
				tsetup_RAD4_ADRCLK_noedge_posedge, tsetup_RAD4_ADRCLK_noedge_posedge,
				thold_RAD4_ADRCLK_noedge_posedge, thold_RAD4_ADRCLK_noedge_posedge,
				REN_ipd = '1', 
				'/', 
				InstancePath & "/R_SAR", 
				TRUE, 
				TRUE, 
				WARNING ); 
 
    END IF; -- Timing Check Section 
 
rd_viol_flag := (Tviol_RAD_stp_hld_0 or Tviol_RAD_stp_hld_1 or Tviol_RAD_stp_hld_2 or Tviol_RAD_stp_hld_3 or Tviol_RAD_stp_hld_4 or Pviol_ADRCLK ); 
 
 
    ------------------------------------------------------------------- 
    -- Functionality Section 
    ------------------------------------------------------------------- 
 
 
if (first) then 
          while( not(endfile(STF)) ) loop 
                readline(STF,readdata) ; 
                read(readdata,tmp_data) ; 
 
  --for T in 0 to 31 loop 
   -- READLINE (STF,readdata); 
   -- Read (readdata,tmp_data); 
    memory_array(T) <= tmp_data; 
    T := T + 1; 
  end loop; 
end if; 
 
 
-- READ CYCLE VIOLATION EFFECT 
 
    if( rd_viol_flag = 'X' or (REN_ipd'EVENT and REN_ipd = '1' and vecX(RD_ADD))) then 
	--output_delay <= 0 ns; 
	data_out <= x_data; 
    elsif 
 
-- VALID MEMORY READ 
 
     (REN_ipd'EVENT and REN_ipd = '1' and not(rd_viol_flag = 'X') and not (vecX(RD_ADD))) then 
	rd_address := vec2int(RD_ADD); 
	data_out <=  memory_array(rd_address); 
    end if; 
 
 
  END PROCESS; 
 
    ------------------------------------------------------------------------------- 
    -- Temporary output signal should get assigned to the output signal. 
    ------------------------------------------------------------------------------- 
 
    --RDATA <= TRANSPORT data_out after output_delay; 

   PROCESS(data_out, ADRCLK_ipd, REN_ipd)

      VARIABLE GLITCH : VitalGlitchDataType;
      VARIABLE RDATA3_1 : std_logic := 'X';
      VARIABLE RDATA2_1 : std_logic := 'X';
      VARIABLE RDATA1_1 : std_logic := 'X';
      VARIABLE RDATA0_1 : std_logic := 'X';

   BEGIN
       RDATA3_1 := VitalBUF(data_out(3));
       RDATA2_1 := VitalBUF(data_out(2));
       RDATA1_1 := VitalBUF(data_out(1));
       RDATA0_1 := VitalBUF(data_out(0));

     VitalPathDelay01 ( RDATA3, GLITCH, "RDATA3", RDATA3_1,
        Paths => (
        0 => ( ADRCLK_ipd'LAST_EVENT, tpd_ADRCLK_RDATA3, TRUE ),
        1 => ( REN_ipd'LAST_EVENT, tpd_REN_RDATA3, TRUE )),
        DefaultDelay=>VitalZeroDelay01,
        Mode=>VitalInertial,
        XON=>TRUE,
        MsgOn=>TRUE,
        MsgSeverity=>WARNING );

     VitalPathDelay01 ( RDATA2, GLITCH, "RDATA2", RDATA2_1,
        Paths => (
        0 => ( ADRCLK_ipd'LAST_EVENT, tpd_ADRCLK_RDATA2, TRUE ),
        1 => ( REN_ipd'LAST_EVENT, tpd_REN_RDATA2, TRUE )),
        DefaultDelay=>VitalZeroDelay01,
        Mode=>VitalInertial,
        XON=>TRUE,
        MsgOn=>TRUE,
        MsgSeverity=>WARNING );

     VitalPathDelay01 ( RDATA1, GLITCH, "RDATA1", RDATA1_1,
        Paths => (
        0 => ( ADRCLK_ipd'LAST_EVENT, tpd_ADRCLK_RDATA1, TRUE ),
        1 => ( REN_ipd'LAST_EVENT, tpd_REN_RDATA1, TRUE )),
        DefaultDelay=>VitalZeroDelay01,
        Mode=>VitalInertial,
        XON=>TRUE,
        MsgOn=>TRUE,
        MsgSeverity=>WARNING );


     VitalPathDelay01 ( RDATA0, GLITCH, "RDATA0", RDATA0_1,
        Paths => (
        0 => ( ADRCLK_ipd'LAST_EVENT, tpd_ADRCLK_RDATA0, TRUE ),
        1 => ( REN_ipd'LAST_EVENT, tpd_REN_RDATA0, TRUE )),
        DefaultDelay=>VitalZeroDelay01,
        Mode=>VitalInertial,
        XON=>TRUE,
        MsgOn=>TRUE,
        MsgSeverity=>WARNING );

END PROCESS;


END VITAL_VF; 
configuration CFG_R_SAR_VITAL of R_SAR is
        for VITAL_VF
        end for;
end CFG_R_SAR_VITAL;
----------------------------------------------------------------------- 
 
