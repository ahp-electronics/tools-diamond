library verilog;
use verilog.vl_types.all;
entity pp_rx_top is
    port(
        rxclk           : in     vl_logic;
        m_rxclk         : in     vl_logic;
        clk             : in     vl_logic;
        rxrst_n         : in     vl_logic;
        m_rxrst_n       : in     vl_logic;
        rst_n           : in     vl_logic;
        rxd_i           : in     vl_logic_vector(9 downto 0);
        rxd_o           : out    vl_logic_vector(11 downto 0);
        mca_rxd_o       : out    vl_logic_vector(10 downto 0);
        mca_rxd_i       : in     vl_logic_vector(11 downto 0);
        ls_sync_status  : out    vl_logic;
        rudi_invalid    : out    vl_logic;
        rudi_idle       : out    vl_logic;
        rudi_config     : out    vl_logic;
        rx_config_reg   : out    vl_logic_vector(15 downto 0);
        xmit            : in     vl_logic_vector(1 downto 0);
        slave           : in     vl_logic;
        cc_re_o         : out    vl_logic;
        cc_we_o         : out    vl_logic;
        cc_re_i         : in     vl_logic;
        cc_we_i         : in     vl_logic;
        mca_en          : in     vl_logic;
        t_detect_dni    : in     vl_logic;
        t_detect_upi    : in     vl_logic;
        t_detect_dno    : out    vl_logic;
        t_detect_upo    : out    vl_logic;
        align_status    : in     vl_logic;
        local_fault     : in     vl_logic_vector(8 downto 0);
        loopback        : in     vl_logic;
        signal_detect   : in     vl_logic;
        enable_cgalign  : in     vl_logic;
        udf_comma_a     : in     vl_logic_vector(9 downto 0);
        udf_comma_b     : in     vl_logic_vector(9 downto 0);
        udf_comma_mask  : in     vl_logic_vector(9 downto 0);
        uc_mode         : in     vl_logic;
        fc_mode         : in     vl_logic;
        rio_mode        : in     vl_logic;
        pcie_mode       : in     vl_logic;
        xge_mode        : in     vl_logic;
        lsm_disable     : in     vl_logic;
        dec_bypass      : in     vl_logic;
        an_enable       : in     vl_logic;
        match1_d        : in     vl_logic_vector(9 downto 0);
        match2_d        : in     vl_logic_vector(9 downto 0);
        match3_d        : in     vl_logic_vector(9 downto 0);
        match4_d        : in     vl_logic_vector(9 downto 0);
        match2_en       : in     vl_logic;
        match4_en       : in     vl_logic;
        min_ipg_cnt     : in     vl_logic_vector(1 downto 0);
        cc_hwm          : in     vl_logic_vector(3 downto 0);
        cc_lwm          : in     vl_logic_vector(3 downto 0);
        pcie_scram_disable: in     vl_logic;
        pcie_scram_select: in     vl_logic;
        cc_overrun      : out    vl_logic;
        cc_underrun     : out    vl_logic;
        scan_mode       : in     vl_logic;
        BISTRUN_A1      : in     vl_logic;
        BISTFC_A1       : in     vl_logic;
        BISTDONE_A1     : out    vl_logic;
        BISTF_A1        : out    vl_logic
    );
end pp_rx_top;
