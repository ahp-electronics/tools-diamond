library verilog;
use verilog.vl_types.all;
entity sbnx16v1mce is
    port(
        A               : in     vl_logic;
        Z               : out    vl_logic
    );
end sbnx16v1mce;
