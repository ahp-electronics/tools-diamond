library verilog;
use verilog.vl_types.all;
entity SYS_TREES is
    port(
        A               : in     vl_logic;
        Y               : out    vl_logic
    );
end SYS_TREES;
