library verilog;
use verilog.vl_types.all;
entity SCLK_TREE is
    port(
        A               : in     vl_logic;
        Z               : out    vl_logic
    );
end SCLK_TREE;
