library verilog;
use verilog.vl_types.all;
entity njtag_fsm is
    generic(
        st_idl          : integer := 0;
        st_dec          : integer := 1;
        st_inf1         : integer := 3;
        st_inf2         : integer := 2;
        st_inf3         : integer := 6;
        st_shf          : integer := 7;
        st_crc          : integer := 5;
        st_dum          : integer := 4
    );
    port(
        njcmd_dec       : out    vl_logic;
        njcmd_inf1      : out    vl_logic;
        njcmd_inf2      : out    vl_logic;
        njcmd_inf3      : out    vl_logic;
        njtag_cmd       : out    vl_logic;
        njtag_infa      : out    vl_logic;
        njshf_dat0      : out    vl_logic;
        njshf_dat       : out    vl_logic;
        njshf_crc       : out    vl_logic;
        njshf_dum       : out    vl_logic;
        njshf_dat_nd    : out    vl_logic;
        nj_frame_end    : out    vl_logic;
        post_dec        : out    vl_logic;
        post_inf1       : out    vl_logic;
        post_inf2       : out    vl_logic;
        post_inf3       : out    vl_logic;
        post_crc        : out    vl_logic;
        fsm_exec_e      : out    vl_logic;
        fsm_exec_f      : out    vl_logic;
        com_shift_en    : out    vl_logic;
        njfsm_hold      : out    vl_logic;
        nj_dsr_shf      : out    vl_logic;
        decom_last_mask : out    vl_logic;
        dum_dat         : out    vl_logic_vector(7 downto 0);
        njtag_slow_response: out    vl_logic;
        njs_halt        : out    vl_logic;
        nj_shf_done     : out    vl_logic;
        nj_last_byte    : out    vl_logic;
        NDUM_DEFAULT    : in     vl_logic_vector(3 downto 0);
        por             : in     vl_logic;
        smclk           : in     vl_logic;
        nj_rst_sync     : in     vl_logic;
        nj_exec_b       : in     vl_logic;
        njport_init     : in     vl_logic;
        njtag_bse_en    : in     vl_logic;
        njtag_slv_en    : in     vl_logic;
        cfg_mstr_busy   : in     vl_logic;
        p_scpu          : in     vl_logic;
        ctrl_srme       : in     vl_logic;
        ctrl_stx_dum    : in     vl_logic_vector(1 downto 0);
        busy_int        : in     vl_logic;
        njtag_data_byte : in     vl_logic_vector(15 downto 0);
        njtag_run       : in     vl_logic;
        njsel_com       : in     vl_logic;
        njsel_dsr       : in     vl_logic;
        cmd_noop        : in     vl_logic;
        nj_cmd_ndata    : in     vl_logic;
        nj_cmd_read     : in     vl_logic;
        nj_cmd_incr     : in     vl_logic;
        nj_cmd_prog     : in     vl_logic;
        nj_cmd_prog_incr: in     vl_logic;
        nj_cmd_read_incr: in     vl_logic;
        nj_cmd_prog_dsr : in     vl_logic;
        nj_cmd_read_dsr : in     vl_logic;
        nj_cmd_read_fslow: in     vl_logic;
        lsc_ebr_read_c  : in     vl_logic;
        lsc_bitstream_burst_c: in     vl_logic;
        lsc_pcs_rw_c    : in     vl_logic;
        lsc_pcs_write_c : in     vl_logic;
        lsc_pcs_read_c  : in     vl_logic;
        sed_cmd_read_incr: in     vl_logic;
        extra_dsr_cnt   : in     vl_logic;
        nj_check_crc_en : in     vl_logic;
        nj_load_op2     : in     vl_logic;
        nj_load_op3     : in     vl_logic;
        njtag_din       : in     vl_logic_vector(7 downto 0);
        nj_operand1     : in     vl_logic_vector(7 downto 0);
        nj_operand2     : in     vl_logic_vector(7 downto 0);
        dsr_cnt_en      : in     vl_logic;
        decompress_njtag_en: in     vl_logic;
        nj_dat_ren      : in     vl_logic;
        nj_dat_wen      : in     vl_logic;
        lsc_sdm         : in     vl_logic;
        finish_bse      : in     vl_logic;
        njburst_inp     : out    vl_logic;
        dec_load        : in     vl_logic
    );
end njtag_fsm;
