library verilog;
use verilog.vl_types.all;
entity efb_pll_sci is
    generic(
        awidth          : integer := 8;
        dwidth          : integer := 8
    );
    port(
        rst_n           : in     vl_logic;
        scan_mode       : in     vl_logic;
        sci_initen      : in     vl_logic_vector(1 downto 0);
        ctrl_tran_ip    : in     vl_logic;
        mc1_sci_part_cfg: in     vl_logic;
        mc1_pll_swap    : in     vl_logic;
        sciclk          : out    vl_logic;
        sciclk_tree     : out    vl_logic;
        wb_clk_i        : in     vl_logic;
        wb_rst_i        : in     vl_logic;
        wb_cyc_i        : in     vl_logic;
        wb_stb_i        : in     vl_logic;
        wb_we_i         : in     vl_logic;
        wb_adr_i        : in     vl_logic_vector;
        wb_dat_i        : in     vl_logic_vector;
        wb_dat_o        : out    vl_logic_vector;
        wb_ack_o        : out    vl_logic;
        cfg_clk_i       : in     vl_logic;
        cfg_rst_i       : in     vl_logic;
        cfg_stb_i       : in     vl_logic;
        cfg_we_i        : in     vl_logic;
        cfg_adr_i       : in     vl_logic_vector;
        cfg_dat_i       : in     vl_logic_vector;
        cfg_dat_o       : out    vl_logic_vector;
        cfg_ack_o       : out    vl_logic;
        pll0_rst_o      : out    vl_logic;
        pll0_stb_o      : out    vl_logic;
        pll0_we_o       : out    vl_logic;
        pll0_adr_o      : out    vl_logic_vector(4 downto 0);
        pll0_dat_o      : out    vl_logic_vector(7 downto 0);
        pll0_dat_i      : in     vl_logic_vector(7 downto 0);
        pll0_ack_i      : in     vl_logic;
        pll1_rst_o      : out    vl_logic;
        pll1_stb_o      : out    vl_logic;
        pll1_we_o       : out    vl_logic;
        pll1_adr_o      : out    vl_logic_vector(4 downto 0);
        pll1_dat_o      : out    vl_logic_vector(7 downto 0);
        pll1_dat_i      : in     vl_logic_vector(7 downto 0);
        pll1_ack_i      : in     vl_logic;
        i2ccr1_1st      : out    vl_logic_vector(7 downto 2);
        i2ccmdr_1st     : out    vl_logic_vector(7 downto 2);
        i2cbr_1st       : out    vl_logic_vector(9 downto 0);
        i2ctxdr_1st     : out    vl_logic_vector(7 downto 0);
        i2ccr1_2nd      : out    vl_logic_vector(7 downto 2);
        i2ccmdr_2nd     : out    vl_logic_vector(7 downto 2);
        i2cbr_2nd       : out    vl_logic_vector(9 downto 0);
        i2ctxdr_2nd     : out    vl_logic_vector(7 downto 0);
        spicr0          : out    vl_logic_vector(7 downto 0);
        spicr1          : out    vl_logic_vector(7 downto 4);
        spicr2          : out    vl_logic_vector(7 downto 0);
        spibr           : out    vl_logic_vector(5 downto 0);
        spicsr          : out    vl_logic_vector(7 downto 0);
        spitxdr         : out    vl_logic_vector(7 downto 0);
        tc_single_shot_mode: out    vl_logic;
        tc_to_reboot_en : out    vl_logic;
        tc_to_reboot_mode: out    vl_logic;
        tc_sclk_sel     : out    vl_logic_vector(2 downto 0);
        tc_cclk_sel     : out    vl_logic_vector(2 downto 0);
        tc_gsrn_dis     : out    vl_logic;
        tc_rstn_ena     : out    vl_logic;
        tc_mode         : out    vl_logic_vector(1 downto 0);
        tc_oc_mode      : out    vl_logic_vector(1 downto 0);
        tc_top_sel      : out    vl_logic;
        tc_ic_ena       : out    vl_logic;
        tc_ovf_ena      : out    vl_logic;
        tc_top_set      : out    vl_logic_vector(15 downto 0);
        tc_ocr_set      : out    vl_logic_vector(15 downto 0);
        tc_cnt_pause    : out    vl_logic;
        tc_cnt_reset    : out    vl_logic;
        tc_oc_force     : out    vl_logic;
        wbccr           : out    vl_logic_vector(7 downto 6);
        wbctxdr         : out    vl_logic_vector(7 downto 0);
        i2csr_1st_sts   : in     vl_logic_vector(7 downto 0);
        i2cgcdr_1st_sts : in     vl_logic_vector(7 downto 0);
        i2crxdr_1st_sts : in     vl_logic_vector(7 downto 0);
        i2csr_2nd_sts   : in     vl_logic_vector(7 downto 0);
        i2cgcdr_2nd_sts : in     vl_logic_vector(7 downto 0);
        i2crxdr_2nd_sts : in     vl_logic_vector(7 downto 0);
        spisr_sts       : in     vl_logic_vector(7 downto 0);
        spirxdr_sts     : in     vl_logic_vector(7 downto 0);
        tc_cnt_sts      : in     vl_logic_vector(15 downto 0);
        tc_top_sts      : in     vl_logic_vector(15 downto 0);
        tc_ocr_sts      : in     vl_logic_vector(15 downto 0);
        tc_icr_sts      : in     vl_logic_vector(15 downto 0);
        tc_ovf_sts      : in     vl_logic;
        tc_ocrf_sts     : in     vl_logic;
        tc_icrf_sts     : in     vl_logic;
        tc_btf_sts      : in     vl_logic;
        wbcsr_sts       : in     vl_logic_vector(7 downto 0);
        wbcrxdr_sts     : in     vl_logic_vector(7 downto 0);
        stb_i2ccr1_1st  : out    vl_logic;
        stb_i2ccmdr_1st : out    vl_logic;
        stb_i2cbr_1st   : out    vl_logic;
        stb_i2ctxdr_1st : out    vl_logic;
        stb_i2cgcdr_1st_sts: out    vl_logic;
        stb_i2crxdr_1st_sts: out    vl_logic;
        stb_i2ccr1_2nd  : out    vl_logic;
        stb_i2ccmdr_2nd : out    vl_logic;
        stb_i2cbr_2nd   : out    vl_logic;
        stb_i2ctxdr_2nd : out    vl_logic;
        stb_i2cgcdr_2nd_sts: out    vl_logic;
        stb_i2crxdr_2nd_sts: out    vl_logic;
        stb_spicr0      : out    vl_logic;
        stb_spicr1      : out    vl_logic;
        stb_spicr2      : out    vl_logic;
        stb_spibr       : out    vl_logic;
        stb_spicsr      : out    vl_logic;
        stb_spitxdr     : out    vl_logic;
        stb_spirxdr_sts : out    vl_logic;
        stb_wbccr       : out    vl_logic;
        stb_wbctxdr     : out    vl_logic;
        stb_wbcrxdr_sts : out    vl_logic;
        i2c_1st_int     : out    vl_logic;
        i2c_2nd_int     : out    vl_logic;
        spi_int         : out    vl_logic;
        timercounter_int: out    vl_logic;
        wbcfg_int       : out    vl_logic;
        passwordThrDetEnable: out    vl_logic;
        accessLockSectorDetEnable: out    vl_logic;
        illegalManuModeDetEnable: out    vl_logic;
        JTAGThrDetEnable: out    vl_logic;
        slaveSPIThrDetEnable: out    vl_logic;
        slaveI2CThrDetEnable: out    vl_logic;
        wishboneThrDetEnable: out    vl_logic
    );
end efb_pll_sci;
