library verilog;
use verilog.vl_types.all;
entity vhiv1mce is
    port(
        Z               : out    vl_logic
    );
end vhiv1mce;
