--
@ER--B$FbsEHo0OR52gR4g-cRRj.jd$R1MHbDO$H0ROQM
R--fN]C8:CsR#//$DMbH0OH$N/lb..jjDjdNl0/NCbbsN#/0D0/HoL/CFM_sdONON/slI_s38PEyf4R

--
-
-
R--1bHlD)CRqIvRHR0E#oHMDqCR7 7)1V1RFssRCRN8NRM8I0sHC-
-RsaNoRC0:kRpO0CMRm-R)RBqd-B
-H
DLssN$CRHC
C;kR#CHCCC38#0_oDFH4O_43ncN;DD
Ck#RCHCC03#8F_Do_HO#MHoCN83D
D;kR#CHCCC38#0_oDFHNO_sEH03DND;H
DLssN$sRFO;Nd
Ck#ROFsNFd3sOONF3lbN;DD
0CMHR0$)_qv)HWR#R
RRCRoMHCsO
R5RRRRRRRRVHNlDR$:#H0sM:oR=MR"F"MC;R
RRRRRRHRI8R0E:MRH0CCos=R:RR(;
RRRRRRRR8N8s8IH0:ERR0HMCsoCRR:=(R;RRRRRR-R-RoLHRFCMkRoEVRFs80CbER
RRRRRRCR8bR0E:MRH0CCos=R:R.R4UR;
RRRRR8RRF_k0sRCo:FRLFNDCM=R:RDVN#RC;RRRR-E-RNF#Rkk0b0CRsoR
RRRRRRHR8MC_soRR:LDFFCRNM:V=RNCD#;RRRR-RR-NRE#NR80HNRM0bkRosC
RRRRRRRR8N8sC_soRR:LDFFCRNM:V=RNCD#RRRRR-R-R8ENRNsC88RN8#sC#CRsoR
RRRRRR;R2
RRRRsbF0
R5RRRRRRRR7amzRRR:FRk0#_08DHFoOC_POs0F58IH04E-RI8FMR0Fj
2;RRRRRRRR7RQhRRR:HRMR#_08DHFoOC_POs0F58IH04E-RI8FMR0Fj
2;RRRRRRRRq)77RRR:HRMR#_08DHFoOC_POs0F58N8s8IH04E-RI8FMR0Fj
2;RRRRRRRRWR RRRR:HRMR#_08DHFoOR;RRRRRRR--I0sHCMRCNCLDRsVFRlsN
RRRRRRRRiBpR:RRRRHMR8#0_oDFHRO;RRRRR-R-RFODOV	RFssRNRl,Ns88,HR8MR
RRRRRRBRmpRiR:MRHR0R#8F_DoRHORRRRR-RR-bRF0DROFRO	VRFs80Fk
RRRRRRRR
2;CRM8CHM00)$Rq)v_W
;
---
-HRwsR#0HDlbCMlC0HN0FlMRkR#0LOCRNCDD8sRNO
Ej-N-
sHOE00COkRsCNEsOjVRFRv)q_R)WHO#
F0M#NRM0M_klODCD#C_8C:bRR0HMCsoCRR:=5C58bR0E-2R4/2d.;RRRRRRRR-R-RFyRVFRsIF#RVBR) Xd.cCRODRD#M8CCCO8
F0M#NRM0M_klODCD#H_I8:CRR0HMCsoCRR:=5H5I8R0E-2R4/;c2RRRRRRRRR-R-RFyRVFRODMkl#VRFR )Bdc.XRDOCDM#RCCC88$
0bFCRkL0_k0#_$RbCHN#Rs$sNRk5MlC_OD_D#8bCCRI8FMR0Fj5,RM_klODCD#H_I8cC*2R+d8MFI0jFR2VRFR8#0_oDFH
O;#MHoNFDRkL0_kR#RRF:RkL0_k0#_$;bCRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-7R.RsNsNF$RVFR8k50RHkMb0FR0RH0s-N#002C#
o#HMRNDF_k0CRMRRRR:#_08DHFoOC_POs0F5lMk_DOCD8#_CRCb8MFI0jFR2R;R-C-RMDNLCV#RF0sRs#H-0CN0#H
#oDMNRCIbjM_CR:RRR8#0_oDFHPO_CFO0sk5MlC_OD_D#8bCCRI8FMR0FjR2;RR--I0sHCMRCNCLD#FRVsNRCOsERFFIRVqR)vCROD
D##MHoNIDRb_C4CRMRR#:R0D8_FOoH_OPC05FsM_klODCD#C_8C8bRF0IMF2Rj;-RR-sRIHR0CCLMNDRC#VRFsCENORIsFRRFV)RqvODCD#H
#oDMNR_HMsRCoR:RRR8#0_oDFHPO_CFO0sH5I8+0EdFR8IFM0R;j2RRRRRRRRRR--k8#CRR0FsHCo#s0CRh7QRH
#oDMNR0Fk_osCR:RRR8#0_oDFHPO_CFO0sH5I8+0EdFR8IFM0R;j2RRRRRRRRRR--k8#CRR0FsHCo#s0CRz7maH
#oDMNR_W )4 tR:RRR8#0_oDFH
O;#MHoNHDRMC_soR4RR#:R0D8_FOoH_OPC05FsI0H8ER+d8MFI0jFR2R;RR#R
HNoMD8RN_osCRRRR:0R#8F_Do_HOP0COFNs58I8sHE80-84RF0IMF2Rj;RRRR-R-RCk#8FR0RosCHC#0s7Rq7#)
HNoMDFRDI8_N8RsR:0R#8F_Do_HOP0COFcs5RI8FMR0FjR2;RRRRRRRRRRRRR-R-R8N8sHRL0H#RM0bkRR0F)RqvODCD#6R5R0LH#CRsJskHC
820C$bRb0l_8N8s$_0bHCR#sRNsRN$5lMk_DOCD8#_CRCb8MFI0jFR2VRFR8#0_oDFHPO_CFO0sgR5RI8FMR0Fj
2;#MHoN0DRlNb_8R8sR0:RlNb_8_8s0C$b;L

CMoH
R
RR-R-RRQVNs88I0H8ERR<6#RN#MHoR''jRR0Fk#MkCL8RH
0#RRRRzR4R:VRHR85N8HsI8R0E=2R4RMoCC0sNCR
RRRRRRFRDI8_N8<sR=jR"j"jjRN&R8C_so25j;R
RRMRC8CRoMNCs0zCR4R;
RzRR.:RRRRHV58N8s8IH0=ERRR.2oCCMsCN0
RRRRRRRRIDF_8N8s=R<Rj"jj&"RR_N8s5Co4FR8IFM0R;j2
RRRR8CMRMoCC0sNC.Rz;R
RRdRzRRR:H5VRNs88I0H8ERR=do2RCsMCN
0CRRRRRRRRD_FINs88RR<=""jjRN&R8C_soR5.8MFI0jFR2R;
RCRRMo8RCsMCNR0Cz
d;RRRRzRcR:VRHR85N8HsI8R0E=2RcRMoCC0sNCR
RRRRRRFRDI8_N8<sR=jR''RR&Ns8_Cdo5RI8FMR0Fj
2;RRRRCRM8oCCMsCN0R;zc
RRRRRz6RH:RVNR58I8sHE80Rc>R2CRoMNCs0RC
RRRRRDRRFNI_8R8s<N=R8C_soR5c8MFI0jFR2R;
RCRRMo8RCsMCNR0Cz
6;
RRRRR--Q5VR8_HMs2CoRosCHC#0sQR7h#RkHRMoB
piRRRRzRnR:VRHRH58MC_soo2RCsMCN
0CRRRRRRRRbOsFCR##5iBp,QR7hL2RCMoH
RRRRRRRRRRRRRHV5iBpR'=R4N'RMB8RpCi'P0CM2ER0CRM
RRRRRRRRRRRRRHRRMC_so=R<Rj5"j"jjR7&RQ;h2
RRRRRRRRRRRR8CMR;HV
RRRRRRRR8CMRFbsO#C#;R
RRMRC8CRoMNCs0zCRnR;
RzRR(:RRRRHV50MFRM8H_osC2CRoMNCs0RC
RRRRRRRRRHRRMC_so=R<Rj5"j"jjR7&RQ;h2
RRRR8CMRMoCC0sNC(Rz;R

RbRRsCFO#5#RB,piR,W R_HMs2CoRoLCHRM
RRRRRHRRVBR5p=iRR''4R8NMRiBp'CCPMR020MEC
RRRRRRRRRRRR_W )4 tRR<=W
 ;RRRRRRRRRRRRHsM_CRo4<H=RMC_soR;
RRRRRCRRMH8RVR;
RCRRMb8RsCFO#
#;
RRRRR--Q5VRNs88_osC2CRso0H#CqsR7R7)kM#HopRBiR
RR4Rz.:RRRRHV58N8sC_soo2RCsMCN
0CRRRRRRRRbOsFCR##5iBp,7Rq7R)2LHCoMR
RRRRRRRRRRVRHRp5BiRR='R4'NRM8B'piCMPC002RE
CMRRRRRRRRRRRRRRRRNs8_C<oR=7Rq7N)58I8sHE80-84RF0IMF2Rj;R
RRRRRRRRRRMRC8VRH;R
RRRRRRMRC8sRbF#OC#R;
RCRRMo8RCsMCNR0Cz;4.
R
RR4RzdRR:H5VRMRF0Ns88_osC2CRoMNCs0RC
RRRRRRRRRNRR8C_so=R<R7q7)85N8HsI8-0E4FR8IFM0R;j2
RRRR8CMRMoCC0sNC4Rzd
;
RRRRzR.nRH:RV8R5F_k0s2CoRMoCC0sNCR
RRRRRRsRbF#OC#mR5B,piR0Fk_osC2CRLo
HMRRRRRRRRRRRRH5VRmiBpR'=R4N'RMm8RB'piCMPC002RE
CMRRRRRRRRRRRRRRRR7amzRR<=F_k0s5CoI0H8ER-48MFI0jFR2R;
RRRRRRRRRCRRMH8RVR;
RRRRRCRRMb8RsCFO#
#;RRRRCRM8oCCMsCN0Rnz.;R

R-RR-CRtMNCs00CRE#CRCODC0FRDo
HORRRRzR4c:FRVsRRHHMMRkOl_C#DD_C8CbFR8IFM0RojRCsMCN
0CRRRR-A-Rk8HDR0FkbRk0CLMND#CRCODC0FRDo
HORRRRRRRR-Q-RVNR58I8sHE80R4>R682RF0M'RCk#RQ1pBCROD
D#RRRRRRRRmn 4RH:RVNR58I8sHE80R4>R6o2RCsMCN
0CRRRRRRRRRRRRRRRRF_k0CHM52=R<R''4RCIEMNR58C_so85N8HsI8-0E4FR8IFM0RR62=2RHR#CDCjR''R;
RRRRRCRRMo8RCsMCNR0Cmn 4;R
RRRRRR-R-RRQV58N8s8IH0>ERRR62qRh758N8s8IH0<ER=6R42#RkCpR1QOBRC#DD
RRRRRRRR4m 6RR:H5VRNs88I0H8ERR=4R62oCCMsCN0
RRRRRRRRRRRRRRRRb0l_8N8s25H58gRF0IMF2RjRR<=h5maOPFM_8#0_oDFHPO_CFO0s,5HR24j2mRX)8RN_osC58N8s8IH04E-RI8FMR0F6
2;RRRRRRRRRRRRRRRR17qh_R46:qR1hj74RsbF0NRlbqR5RR=>0_lbNs8855H2jR2,A>R=Rb0l_8N8s25H5,42R=BR>lR0b8_N8Hs5225.,RR7=0>RlNb_858sHd252R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR =0>RlNb_858sHc252w,RRR=>0_lbNs8855H26R2,t>R=Rb0l_8N8s25H5,n2R=]R>lR0b8_N8Hs5225(,RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRQ=0>RlNb_858sHU252K,RRR=>0_lbNs8855H2gR2,Z>R=R0Fk_5CMH;22
RRRRRRRR8CMRMoCC0sNC Rm4
6;RRRRRRRRmc 4RH:RVNR58I8sHE80R4=Rco2RCsMCN
0CRRRRRRRRRRRRRRRR0_lbNs8855H2UFR8IFM0RRj2<h=RmOa5F_MP#_08DHFoOC_POs0F5RH,gR22XRm)Ns8_CNo58I8sHE80-84RF0IMF2R6;R
RRRRRRRRRRRRRRqR1h47_cRR:17qh4bjRFRs0lRNb5=qR>lR0b8_N8Hs5225j,RRA=0>RlNb_858sH4252B,RRR=>0_lbNs8855H2.R2,7>R=Rb0l_8N8s25H5,d2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR >R=Rb0l_8N8s25H5,c2R=wR>lR0b8_N8Hs52256,RRt=0>RlNb_858sHn252],RRR=>0_lbNs8855H2(R2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRQ>R=Rb0l_8N8s25H5,U2R=KR>4R''Z,RRR=>F_k0CHM52
2;RRRRRRRRCRM8oCCMsCN0R4m cR;
RRRRRmRR R4d:VRHR85N8HsI8R0E=dR42CRoMNCs0RC
RRRRRRRRRRRRR0RRlNb_858sH(25RI8FMR0Fj<2R=mRhaF5OM#P_0D8_FOoH_OPC05FsHU,R2X2RmN)R8C_so85N8HsI8-0E4FR8IFM0R;62
RRRRRRRRRRRRRRRRh1q7d_4R1:RqUh7RFRbsl0RN5bRq>R=Rb0l_8N8s25H5,j2R=AR>lR0b8_N8Hs52254,RRB=0>RlNb_858sH.2527,RRR=>0_lbNs8855H2d
2,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR RRRR=>0_lbNs8855H2cR2,w>R=Rb0l_8N8s25H5,62R=tR>lR0b8_N8Hs5225n,RR]=0>RlNb_858sH(252
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRZRRRR=>F_k0CHM52
2;RRRRRRRRCRM8oCCMsCN0R4m dR;
RRRRRmRR R4.:VRHR85N8HsI8R0E=.R42CRoMNCs0RC
RRRRRRRRRRRRR0RRlNb_858sHn25RI8FMR0Fj<2R=mRhaF5OM#P_0D8_FOoH_OPC05FsH(,R2X2RmN)R8C_so85N8HsI8-0E4FR8IFM0R;62
RRRRRRRRRRRRRRRRh1q7._4R1:RqUh7RFRbsl0RN5bRq>R=Rb0l_8N8s25H5,j2R=AR>lR0b8_N8Hs52254,RRB=0>RlNb_858sH.2527,RRR=>0_lbNs8855H2d
2,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR RRRR=>0_lbNs8855H2cR2,w>R=Rb0l_8N8s25H5,62R=tR>lR0b8_N8Hs5225n,RR]='>R4R',
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRZ>R=R0Fk_5CMH;22
RRRRRRRR8CMRMoCC0sNC Rm4
.;RRRRRRRRm4 4RH:RVNR58I8sHE80R4=R4o2RCsMCN
0CRRRRRRRRRRRRRRRR0_lbNs8855H26FR8IFM0RRj2<h=RmOa5F_MP#_08DHFoOC_POs0F5RH,nR22XRm)Ns8_CNo58I8sHE80-84RF0IMF2R6;R
RRRRRRRRRRRRRRqR1h47_4RR:17qhnbRRFRs0lRNb5=qR>lR0b8_N8Hs5225j,RRA=0>RlNb_858sH4252B,RRR=>0_lbNs8855H2.R2,7>R=Rb0l_8N8s25H5,d2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR >R=Rb0l_8N8s25H5,c2R=wR>lR0b8_N8Hs52256,RRZ=F>RkC0_M25H2R;
RRRRRCRRMo8RCsMCNR0Cm4 4;R
RRRRRR Rm4:jRRRHV58N8s8IH0=ERR24jRMoCC0sNCR
RRRRRRRRRRRRRRlR0b8_N8Hs52R5c8MFI0jFR2=R<Rahm5MOFP0_#8F_Do_HOP0COFHs5,2R62mRX)8RN_osC58N8s8IH04E-RI8FMR0F6
2;RRRRRRRRRRRRRRRR17qh_R4j:qR1hR7nRsbF0NRlbqR5RR=>0_lbNs8855H2jR2,A>R=Rb0l_8N8s25H5,42R=BR>lR0b8_N8Hs5225.,RR7=0>RlNb_858sHd252R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR =0>RlNb_858sHc252w,RRR=>',4'R=ZR>kRF0M_C52H2;R
RRRRRRMRC8CRoMNCs0mCR ;4j
RRRRRRRRgm RRR:H5VRNs88I0H8ERR=go2RCsMCN
0CRRRRRRRRRRRRRRRR0_lbNs8855H2dFR8IFM0RRj2<h=RmOa5F_MP#_08DHFoOC_POs0F5RH,cR22XRm)Ns8_CNo58I8sHE80-84RF0IMF2R6;R
RRRRRRRRRRRRRRqR1hg7_R1:Rqch7RbRRFRs0lRNb5=qR>lR0b8_N8Hs5225j,RRA=0>RlNb_858sH4252B,RRR=>0_lbNs8855H2.R2,7>R=Rb0l_8N8s25H5,d2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRZ>R=R0Fk_5CMH;22
RRRRRRRR8CMRMoCC0sNC RmgR;
RRRRRmRR RUR:VRHR85N8HsI8R0E=2RURMoCC0sNCR
RRRRRRRRRRRRRRlR0b8_N8Hs52R5.8MFI0jFR2=R<Rahm5MOFP0_#8F_Do_HOP0COFHs5,2Rd2mRX)8RN_osC58N8s8IH04E-RI8FMR0F6
2;RRRRRRRRRRRRRRRR17qh_:URRh1q7RcRRsbF0NRlbqR5RR=>0_lbNs8855H2jR2,A>R=Rb0l_8N8s25H5,42R=BR>lR0b8_N8Hs5225.,RR7='>R4
',RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRZRRRR=>F_k0CHM52
2;RRRRRRRRCRM8oCCMsCN0RUm ;R
RRRRRR Rm(:RRRRHV58N8s8IH0=ERRR(2oCCMsCN0
RRRRRRRRRRRRRRRRb0l_8N8s25H584RF0IMF2RjRR<=h5maOPFM_8#0_oDFHPO_CFO0s,5HR2.2R)XmR_N8s5CoNs88I0H8ER-48MFI06FR2R;
RRRRRRRRRRRRR1RRq_h7(RR:17qh.RRRb0FsRblNRR5q=0>RlNb_858sHj252A,RRR=>0_lbNs8855H24R2,Z>R=R0Fk_5CMH;22
RRRRRRRR8CMRMoCC0sNC Rm(R;
RRRRRmRR RnR:VRHR85N8HsI8R0E=2RnRMoCC0sNCR
RRRRRRRRRRRRRRkRF0M_C5RH2<'=R4I'RERCM5_N8s5Co6=2RRMOFP0_#8F_Do_HOP0COFHs5,542jR22CCD#R''j;R
RRRRRRMRC8CRoMNCs0mCR 
n;RRRR-Q-RVNR58I8sHE80RR<=6M2RFkRF00bkRNCMLRDC#CCDOD0RFOoHRCMC8RC8/NRlbHR8s0COD0$RFqR)vR'#Ns88CR##DCHM#R
RRRRRR Rm6RR:H5VRNs88I0H8E=R<RR62oCCMsCN0
RRRRRRRRRRRRRRRR0Fk_5CMH<2R=4R''R;
RRRRRCRRMo8RCsMCNR0Cm; 6
R
RR-R-RRQV58N8s8IH0>ERRRg2kR#CWju RR0F8FCO8NCR8C8s#L#RHR0#nER0soFkERRgNRM8W4u RR0F8FCO8LCRHR0#4+jR
RRRRRRRR4W jRR:H5VRNs88I0H8ERR>go2RCsMCN
0CRRRRRRRRRRRRRRRRIjbC_5CMH<2R=4R''ERIC5MRNs8_CUo5RI8FMR0F6=2RRMOFP0_#8F_Do_HOP0COFHs5,2.j58dRF0IMF2Rj2DRC#'CRj
';RRRRRRRRRRRRRRRRI4bC_5CMH<2R=4R''ERIC5MRNs8_CNo58I8sHE80-84RF0IMF2RgRO=RF_MP#_08DHFoOC_POs0F5.H,jN258I8sHE80-8nRF0IMF2Rc2DRC#'CRj
';RRRRRRRRRRRRCRM8oCCMsCN0R4W jR;
R-RR-VRQR85N8HsI8R0E=RRUFgsR2#RkCuRW 0jRFCR8OCF8R8N8s#C#R0LH#RRn0FEskRoEgR
RRRRRR RWg:RRRRHV585N8HsI8R0E=2RURRm)58N8s8IH0=ERR2g2RMoCC0sNCR
RRRRRRRRRRRRRRbRICCj_M25HRR<='R4'IMECR85N_osC58N8s8IH04E-RI8FMR0F6=2RRRH2CCD#R''j;R
RRRRRRRRRRRRRRbRICC4_M25HRR<=';4'
RRRRRRRRRRRR8CMRMoCC0sNC RWgR;
R-RR-VRQR85N8HsI8R0E=2R(RCk#R WujFR0RO8CFR8C0RECnR0ENs88CR##LRH0&uRW 04RFCR8OCF8RC0ERE(0R8N8s#C#R0LH
RRRRRRRR(W RRR:H5VRNs88I0H8ERR=(o2RCsMCN
0CRRRRRRRRRRRRRRRRIjbC_5CMH<2R=4R''ERIC5MRNs8_C6o52RR=OPFM_8#0_oDFHPO_CFO0s,5H.j252C2RDR#C';j'
RRRRRRRRRRRRRRRRCIb4M_C5RH2<'=R4I'RERCM5_N8s5Con=2RRMOFP0_#8F_Do_HOP0COFHs5,5.24R22CCD#R''j;R
RRRRRRMRC8CRoMNCs0WCR 
(;RRRR-Q-RVNR58I8sHE80Rn=R2#RkCuRW 0jRFCR8OCF8RC0EREn0R8N8s#C#R0LH
RRRRRRRRnW RRR:H5VRNs88I0H8ERR=no2RCsMCN
0CRRRRRRRRRRRRRRRRIjbC_5CMH<2R=4R''ERIC5MRNs8_C6o52RR=OPFM_8#0_oDFHPO_CFO0s,5H4j252C2RDR#C';j'
RRRRRRRRRRRRRRRRCIb4M_C5RH2<'=R4
';RRRRRRRRCRM8oCCMsCN0RnW ;R
RR-R-RRQV58N8s8IH0<ER=2R6RRMFI0sHCMRCNCLDRD#CCRO0DHFoOCRMC88C
RRRRRRRR6W RRR:H5VRNs88I0H8E=R<RR62oCCMsCN0
RRRRRRRRRRRRRRRRCIbjM_C5RH2<'=R4
';RRRRRRRRRRRRRRRRI4bC_5CMH<2R=4R''R;
RRRRRCRRMo8RCsMCNR0CW; 6
R
RRMRC8CRoMNCs0zCR4
c;
RRRR6z.RH:RVMR5F80RF_k0s2CoRMoCC0sNCR
RRRRRR4Rz(R4:bOsFCR##5_W )4 t,MRH_osC4F,Rks0_C
o2RRRRRRRRLHCoMR
RRRRRRRRRRVRHR 5W_t) 4RR='24'RC0EMR
RRRRRRRRRRRRRRmR7z<aR=MRH_osC4H5I8-0E4FR8IFM0R;j2
RRRRRRRRRRRR#CDCR
RRRRRRRRRRRRRRmR7z<aR=kRF0C_soH5I8-0E4FR8IFM0R;j2
RRRRRRRRRRRR8CMR;HV
RRRRRRRR8CMRFbsO#C#R(z44R;
RCRRMo8RCsMCNR0Cz;.6
R
RR-R-RMtCC0sNCER0CqR)vCRODRD#IEH0RH0s-N#00
C#RRRRzR46:FRVsRRHHMMRkOl_C#DD_C8CbFR8IFM0RojRCsMCN
0CRRRRRRRRzR4(:FRVsRR[HMMRkOl_C#DD_8IHCFR8IFM0RojRCsMCN
0CRRRRRRRRRRRRzv)q:BR) Xd.cRR
RRRRRRRRRRRRRbRRFRs0lRNb5j7QRR=>HsM_C5o5[2*c27,RQ=4R>MRH_osC5*5[c42+27,RQ=.R>MRH_osC5*5[c.2+27,RQ=dR>MRH_osC5*5[cd2+2R,
RRRRRRRRRRRRRRRRRRRRRRRRRjq7RR=>D_FINs885,j2R4q7RR=>D_FINs885,42R.q7RR=>D_FINs885,.2Rdq7RR=>D_FINs885,d2Rcq7RR=>D_FINs885,c2
R--RRRRRRRRRRRRRRRRRRRRRRRRR W)h>R=R,W R Wuj>R=RCIbjM_C5,H2R Wu4>R=RCIb4M_C5,H2RRBi=h>RmBaRpRi,
RRRRRRRRRRRRRRRRRRRRRRRRWRR)R h=W>R W,RuR j=I>Rb_CjCHM52W,RuR 4=I>Rb_C4CHM52B,Ri>R=RiBp,1Rt)>R=R''4,RR
RRRRRRRRRRRRRRRRRRRRRRRRRj7mRR=>F_k0L5k#H[,5*2c2,mR74>R=R0Fk_#Lk55H,[2*c+,42R.7mRR=>F_k0L5k#H[,5*+c2.R2,7Rmd=F>RkL0_kH#5,*5[cd2+2
2;RRRRRRRRRRRRRRRRF_k0s5Co5c[*2<2R=kRF0k_L#,5H5c[*2I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co5c[*22+4RR<=F_k0L5k#H[,5*+c24I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co5c[*22+.RR<=F_k0L5k#H[,5*+c2.I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co5c[*22+dRR<=F_k0L5k#H[,5*+c2dI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRCRM8oCCMsCN0R(z4;R
RRRRRRMRC8CRoMNCs0zCR4
6;
R--RUz.RH:RV8R5F_k0s2CoRMoCC0sNC-
-RRRRRRRRzR4n:FRVsRRHHMMRkOl_C#DD_C8CbFR8IFM0RojRCsMCN
0C-R-RRRRRR4RzURR:VRFs[MRHRlMk_DOCDI#_HR8C8MFI0jFRRMoCC0sNC-
-RRRRRRRRRRRRzv)q:BR) Xd.c-R
-RRRRRRRRRRRRRRRRsbF0NRlb7R5Q=jR>MRH_osC5*5[c,22R47QRR=>HsM_C5o5[2*c+,42R.7QRR=>HsM_C5o5[2*c+,.2Rd7QRR=>HsM_C5o5[2*c+,d2
R--RRRRRRRRRRRRRRRRRRRRRRRRRjq7RR=>D_FINs885,j2R4q7RR=>D_FINs885,42R.q7RR=>D_FINs885,.2Rdq7RR=>D_FINs885,d2Rcq7RR=>D_FINs885,c2
R--RRRRRRRRRRRRRRRRRRRRRRRRR W)h>R=R,W R Wuj>R=RCIbjM_C5,H2R Wu4>R=RCIb4M_C5,H2RRBi=h>RmBaRpRi,
R--RRRRRRRRRRRRRRRRRRRRRRRRRmT7j>R=R0Fk_#Lk55H,[2*c2T,R7Rm4=F>RkL0_kH#5,*5[c42+2T,R7Rm.=F>RkL0_kH#5,*5[c.2+2T,R7Rmd=F>RkL0_kH#5,*5[cd2+2
2;-R-RRRRRRRRRRRRRRkRF0C_so[55*2c2RR<=F_k0L5k#H[,5*2c2RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;-
-RRRRRRRRRRRRRRRRF_k0s5Co5c[*22+4RR<=F_k0L5k#H[,5*+c24I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';-R-RRRRRRRRRRRRRRkRF0C_so[55*+c2.<2R=kRF0k_L#,5H5c[*22+.RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;-
-RRRRRRRRRRRRRRRRF_k0s5Co5c[*22+dRR<=F_k0L5k#H[,5*+c2dI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';-R-RRRRRRRRRRMRC8CRoMNCs0zCR4
U;-R-RRRRRR8CMRMoCC0sNC4Rzn-;
-RRRR8CMRMoCC0sNC.RzU
;
-R-RRRRRk:URRRHV5k8F0C_soo2RCsMCN
0C-R-RRRRRRRRR7amzRR<=F_k0s5CoI0H8ER-48MFI0jFR2-;
-CRRMo8RCsMCNR0Ck
U;RRRRRRRRRRRRRRRRRM
C8sRNO0EHCkO0sNCRsjOE;



