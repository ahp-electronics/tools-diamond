library verilog;
use verilog.vl_types.all;
entity config_jtag is
    port(
        pll_set         : in     vl_logic_vector(7 downto 0);
        pll_set2        : in     vl_logic_vector(5 downto 0);
        wake_period     : in     vl_logic_vector(2 downto 0);
        done_phase      : in     vl_logic_vector(3 downto 0);
        goe_phase       : in     vl_logic_vector(2 downto 0);
        gwd_phase       : in     vl_logic_vector(2 downto 0);
        gsr_phase       : in     vl_logic_vector(2 downto 0);
        syn_ext_done    : in     vl_logic;
        prog_128        : in     vl_logic;
        idcode          : in     vl_logic_vector(31 downto 0);
        clear_finish    : in     vl_logic;
        start           : in     vl_logic;
        operation       : in     vl_logic;
        preamble        : in     vl_logic;
        exit_abort      : in     vl_logic;
        illegal_rd      : in     vl_logic;
        por             : in     vl_logic;
        tms             : in     vl_logic;
        tck             : in     vl_logic;
        tdi             : in     vl_logic;
        asrout_0        : in     vl_logic;
        dsrout_0        : in     vl_logic;
        bsout_0         : in     vl_logic;
        cmd_ld_ucode    : in     vl_logic;
        cmd_rd_ucode    : in     vl_logic;
        cmd_prgm_done_r : in     vl_logic;
        cmd_prgm_done_comp: in     vl_logic;
        cmd_prgm_sec    : in     vl_logic;
        cmd_clear_all_r : in     vl_logic;
        cmd_ld_ctrl0    : in     vl_logic;
        cmd_rd_ctrl0    : in     vl_logic;
        crc_err         : in     vl_logic;
        id_fail_r       : in     vl_logic;
        non_jtag_config : in     vl_logic;
        read_back       : in     vl_logic;
        cmd_bypass      : in     vl_logic;
        cmd_flow_thru   : in     vl_logic;
        program         : in     vl_logic;
        mux_clk         : in     vl_logic;
        wakeup_clk      : in     vl_logic;
        cmd_ctrl0_r     : in     vl_logic_vector(31 downto 0);
        cmd_ucode_r     : in     vl_logic_vector(31 downto 0);
        cmd_crc         : in     vl_logic_vector(15 downto 0);
        er1out          : in     vl_logic;
        er2out          : in     vl_logic;
        break_chain     : in     vl_logic;
        clear_memory    : in     vl_logic;
        pll_lock        : in     vl_logic_vector(7 downto 0);
        ext_done        : in     vl_logic;
        cmd_bypass_en   : in     vl_logic;
        pcm             : in     vl_logic;
        serial          : in     vl_logic;
        forcearch       : in     vl_logic;
        pll_lock2       : in     vl_logic_vector(5 downto 0);
        spi_sel         : out    vl_logic_vector(2 downto 0);
        isc_inst_tri    : out    vl_logic;
        async_rst       : out    vl_logic;
        mclk_en_r       : out    vl_logic;
        jtag_active     : out    vl_logic;
        mfgen           : out    vl_logic;
        edit_mod        : out    vl_logic;
        decomp_en       : out    vl_logic;
        auto_clear      : out    vl_logic;
        mck_freq_switch : out    vl_logic;
        progen          : out    vl_logic;
        jtag_data       : out    vl_logic;
        jtag_addr       : out    vl_logic;
        tdo_out         : out    vl_logic;
        tdo_en          : out    vl_logic;
        reg_rd_bus      : out    vl_logic_vector(31 downto 0);
        done_pupb       : out    vl_logic;
        security        : out    vl_logic;
        freq_sel        : out    vl_logic_vector(5 downto 0);
        freq_div        : out    vl_logic_vector(5 downto 0);
        overload        : out    vl_logic_vector(1 downto 0);
        glb_reg_rd      : out    vl_logic;
        init_r          : out    vl_logic;
        nonjtag_cfg_r   : out    vl_logic;
        read_back_r     : out    vl_logic;
        error           : out    vl_logic;
        rst_addr_o      : out    vl_logic;
        rti             : out    vl_logic;
        goe_high_r      : out    vl_logic;
        gwd_high_r      : out    vl_logic;
        gsr_high_r      : out    vl_logic;
        done_high_all   : out    vl_logic;
        exit_start_dly  : out    vl_logic;
        selasr          : out    vl_logic;
        seldsr          : out    vl_logic;
        ipa_o           : out    vl_logic;
        ipb_o           : out    vl_logic;
        iptesta_o       : out    vl_logic;
        iptestb_o       : out    vl_logic;
        erase_o         : out    vl_logic;
        prog_inc_rti_o  : out    vl_logic;
        vfy_incr_rti_o  : out    vl_logic;
        rst_crc_o       : out    vl_logic;
        bsmode1         : out    vl_logic;
        bsmode2         : out    vl_logic;
        bsmode3         : out    vl_logic;
        burst_o         : out    vl_logic;
        wakeup_minus_r  : out    vl_logic;
        wakeup_minus    : out    vl_logic;
        jtag_unprogram  : out    vl_logic;
        jtag_unprogram_dly: out    vl_logic;
        jtag_functional : out    vl_logic;
        shiftdr         : out    vl_logic;
        burst_clear     : out    vl_logic;
        upir            : out    vl_logic;
        capdr           : out    vl_logic;
        updr            : out    vl_logic;
        seldr           : out    vl_logic;
        selir           : out    vl_logic;
        tlreset         : out    vl_logic;
        nonjtag_active  : out    vl_logic;
        done_reg        : out    vl_logic;
        extest          : out    vl_logic;
        sample          : out    vl_logic;
        tdi_bscan       : out    vl_logic;
        selbsr          : out    vl_logic;
        edit_xread      : out    vl_logic;
        test_cntls      : out    vl_logic_vector(55 downto 0);
        init            : out    vl_logic;
        refresh_o       : out    vl_logic
    );
end config_jtag;
