library verilog;
use verilog.vl_types.all;
entity ctr_cntl is
    port(
        HWRITE          : out    vl_logic;
        HWDATA          : out    vl_logic_vector(35 downto 0);
        HSIZE           : out    vl_logic_vector(1 downto 0);
        HRDATA          : out    vl_logic_vector(35 downto 0);
        HGRANT_MPI      : out    vl_logic;
        HGRANT_FPSC     : out    vl_logic;
        HGRANT_FPGA     : out    vl_logic;
        HGRANT_CFG      : out    vl_logic;
        HADDR           : out    vl_logic_vector(17 downto 0);
        HMASTER         : out    vl_logic_vector(3 downto 0);
        HREADY          : out    vl_logic;
        HTRANS          : out    vl_logic_vector(1 downto 0);
        HRESP           : out    vl_logic_vector(1 downto 0);
        HSEL_FPGA       : out    vl_logic;
        HSEL_LFPSC      : out    vl_logic;
        HSEL_RAMT       : out    vl_logic;
        HSEL_RFPSC      : out    vl_logic;
        HSEL_SBC        : out    vl_logic;
        HBURST          : out    vl_logic;
        RASB_SLAVE_ENABLE: in     vl_logic;
        PRIORITY_MPI    : in     vl_logic_vector(1 downto 0);
        PRIORITY_FPSC   : in     vl_logic_vector(1 downto 0);
        PRIORITY_FPGA   : in     vl_logic_vector(1 downto 0);
        PAD_DONE        : in     vl_logic;
        LOCK_USER       : in     vl_logic;
        LOCK_MPI        : in     vl_logic;
        LOCK_FPSC       : in     vl_logic;
        LASB_SLAVE_ENABLE: in     vl_logic;
        HWRITE_MPI      : in     vl_logic;
        HWRITE_FPSC     : in     vl_logic;
        HWRITE_FPGA     : in     vl_logic;
        HWRITE_CFG      : in     vl_logic;
        HWDATA_MPI      : in     vl_logic_vector(35 downto 0);
        HWDATA_FPSC     : in     vl_logic_vector(35 downto 0);
        HWDATA_FPGA     : in     vl_logic_vector(35 downto 0);
        HWDATA_CFG      : in     vl_logic_vector(35 downto 0);
        HTRANS_MPI      : in     vl_logic_vector(1 downto 0);
        HTRANS_FPSC     : in     vl_logic_vector(1 downto 0);
        HTRANS_FPGA     : in     vl_logic_vector(1 downto 0);
        HTRANS_CFG      : in     vl_logic_vector(1 downto 0);
        HSIZE_MPI       : in     vl_logic_vector(1 downto 0);
        HSIZE_FPSC      : in     vl_logic_vector(1 downto 0);
        HSIZE_FPGA      : in     vl_logic_vector(1 downto 0);
        HSIZE_CFG       : in     vl_logic_vector(1 downto 0);
        HRESP_SBC       : in     vl_logic_vector(1 downto 0);
        HRESP_RFPSC     : in     vl_logic_vector(1 downto 0);
        HRESP_RAMT      : in     vl_logic_vector(1 downto 0);
        HRESP_LFPSC     : in     vl_logic_vector(1 downto 0);
        HRESP_FPGA      : in     vl_logic_vector(1 downto 0);
        HRESET_N        : in     vl_logic;
        HREADY_SBC      : in     vl_logic;
        HREADY_RFPSC    : in     vl_logic;
        HREADY_RAMT     : in     vl_logic;
        HREADY_LFPSC    : in     vl_logic;
        HREADY_FPGA     : in     vl_logic;
        HRDATA_SBC      : in     vl_logic_vector(35 downto 0);
        HRDATA_RFPSC    : in     vl_logic_vector(35 downto 0);
        HRDATA_LFPSC    : in     vl_logic_vector(35 downto 0);
        HRDATA_FPGA     : in     vl_logic_vector(35 downto 0);
        HLOCK_MPI       : in     vl_logic;
        HLOCK_FPSC      : in     vl_logic;
        HLOCK_FPGA      : in     vl_logic;
        HLOCK_CFG       : in     vl_logic;
        HCLK_SWITCH     : in     vl_logic;
        HCLK            : in     vl_logic;
        HBUSREQ_MPI     : in     vl_logic;
        HBUSREQ_FPSC    : in     vl_logic;
        HBUSREQ_FPGA    : in     vl_logic;
        HBUSREQ_CFG     : in     vl_logic;
        HADDR_MPI       : in     vl_logic_vector(17 downto 0);
        HADDR_FPSC      : in     vl_logic_vector(17 downto 0);
        HADDR_FPGA      : in     vl_logic_vector(17 downto 0);
        HADDR_CFG       : in     vl_logic_vector(17 downto 0);
        Timeout_Index1  : in     vl_logic_vector(3 downto 0);
        Timeout_Index2  : in     vl_logic_vector(3 downto 0);
        HBURST_CFG      : in     vl_logic;
        HBURST_FPGA     : in     vl_logic;
        HBURST_FPSC     : in     vl_logic;
        HBURST_MPI      : in     vl_logic
    );
end ctr_cntl;
