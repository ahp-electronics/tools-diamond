------------------------------------------------------------------------
@E
---a-RERH#VCHDR#ENRR0FL#CREbHbCC8RM$Osb80C!
!!-a-RERH#VCHDRF#EkRD8MCCPsCRLRH#Eb8bCRRHMs8CNNCLDRsVFl!!!

---a-RERH#P#CsHRFMF0VREvCRq_a]BumvpR Xb	NONRoCH-#
-bR1CVOHH0ORF$R1MHbDVN$RMH8R#FRM0#RkNCLDRsVFRl#Hk0DNH
FM-B-RFsb$H0oER25ORg4gc1,R$DMbH0OH$Q,RMRO3qRDDsEHo0s#RCs#CP
C8---
-ERaC>R=RCFbsFN0s#RHRCk#8FR0RC#bO$HVRLNRk0HDRRHMHDlbCMlC0HN0F
MR-V-RFNsRRb0$CsRFRMVkOF0HM-3
--
-RCaER8FsCFsRVkRVMHO0FRM#NRM88DCON0sNH#FMRRH#MRF0HM8C0NHODFR0RC0E
R--FosHHDMNRsPC#MHFRsVFRO#Ck0sH$CRsNM#F#-3
--
-RCf]Ns8C:/R/#b$MDHHO0O$/F.lbjj.jdM#$bO./FHlbD#Cs/8PEDE/P8N/l0OE_FDlbCPG3E48yR-f
--
-RswFRswk0sECR#8CObsH0MHFR08CN#HD,DRbCCN#RFDF	0RNRlOFl0CM#CRLD:FI
-------------------------------------------------------------------------
-
R--B$FbsEHo0gR4gLnR$ RQ R 3qRDDsEHo0s#RCs#CP3C8

---a-RERH##sFkOVCRHRDCHN#RM#RC#0CMHRNDb0NsRRFVQ   R810R(4jn-3.4ngg, RQ 1 R08NMNRs8
R--ep]7R0vNENCl0NHODNRuOo	NCR#3a#EHRk#FsROCVCHDR$lNR0MFRRLCOHFbCR8,#8FD,sRFR-
-ROHMDCk88HRI0#ERFIV0NRsC00ENRRH##8FDR0IHE0FkRHIs0M0CRsbCl#H#HRFMVlsFRC0ER Q  -
-RN10Ms8N87#RCsbN0MlC0a3RERH##sFkOVCRHRDClRN$LkCR#RC80HFRlCbDl0CMRH0E#0R#NNM8s
8R-N-RMl8RNL$RCHR8#H0sLCk08MRHRlOFbCHD8FRVsHlRMMRN$NRlMsMCRR#FDoFMRRN#0REC
R--ObFlH8DCRsVFlFR8CM#RFN0RDIDFRs8HCRO08FCOlDbHNF0HMVRFRC0ERHFsoNHMDFR#kCsORDVHC-3
-ERaH##RFOksCHRVDlCRNL$RCFROb8HCRsVFR8HMH8PHkRNDkR#CLIC0CRCMDCHOM8#CRCk#sR#3
R--a#EHRk#FsROCVCHDRRH#bPsFH88CRRFMNqMR11RQR#LNHR#3aRECQ   R#8HOHDNlq#Rh
YR-W-Rqq))hRaY )Xu R11mQ)RvQup Q7RhzBp7tQhRYqhR)Wq)aqhYwRmR)v Bh]qaQqApYQaR-
-R7qhRawQh1 1R)wmR z1R)wmRuqRqQ)aBqzp)zRu)1um a3REkCR#RCsF0VRE#CRFOksC-R
-HRVD#CREDNDR8HMCHlMVN$RME8RFRD8Q   RsENl#DC#sRVFNlRM8$RNolNCF#RsHRDNDLHHR0$
R--N#sHHRMoFRk0F0VREkCR#0CRECCsF
V3---
-HRa0:DCRRRRR1RR08NMNRs8ep]7R0vNENCl0NHODNRuOo	NC5#RQ   R810R(4jn-3.4ngg,-
-RRRRRRRRRRRRRqRvaB]_mpvu 
X2---
-HRpLssN$R:RRaRRERH#b	NONRoC#DENDCRLRlOFbCHD8MRH0NFRRLDHs$Ns
R--RRRRRRRRRRRRRl#$LHFDODND$NRMlRC8Q   3-
-
R--7CCPDCFbsR#:R Q  qR71eBR]R7pvEN0C0lNHDONROuN	CNo#FRWsM	HosRtF
kb---
-kRus#bFCR:RRaRRERH#b	NONRoC8HCVMRC#N0R#NNM8sV8RF8sRCo#HM#CsRR0FkR#CH-M
-RRRRRRRRRRRR8RRCs#OHMLHo]Re7lpRFD8C#ER0Nl0RNR	CkR#CFOVRFFllMmRBv upX-
-RRRRRRRRRRRRRFROMN#0MR0#NRM8OlFlFBMRmpvu lXRNC0ElHN0ORNDVOkM0MHF#MRN8-
-RRRRRRRRRRRRRbRFC0sNF3s#

---p-RH0lHNF0HMR:RaRECPkNDCo#RCsMCN80CRRL$0RECVOkM0MHF#MRHRH0E#NRbOo	NCNRl$-
-RRRRRRRRRRRRRNRPsV$RsRFlb0DNVlFsRR0Fb0DNVlFs,MRN8ER0CsRbC#OHHRFMFsVRCD#k0-#
-RRRRRRRRRRRRHRR#MRFDo$RkNNsMC0C8FR0RRLC0REClHHMlRklskCJH8sCRRL$Q   R810R(4jn--
-RRRRRRRRRRRR4RRg3gd

---h-RF#0C:-
-RRRRRRRRRRRRRFRhRO8CDNNs0MHF#sRFRV8CH0MHH#FMRN#EDLDRCMRHO8DkCH8RMF,Rs-
-RRRRRRRRRRRRRGRCO8DkCV8Rs,FlRH0E#NRbOo	NC-3
-RRRRRRRRRRRRaRRE"CRb	NONRoC8DCON0sNH"FMRV8CH#MCRC0ERb0$CR#,#0kL$#bC,MRN8-
-RRRRRRRRRRRRRCR8OsDNNF0HMF#RVqRvaB]_mpvu 
X3-R-RRRRRRRRRRRRRaREC#M0N88NsR0lNENCl0NHODCR8VHHM0MHFR8NMRMOFP0CMHNFMDCRlNMMHo-
-RRRRRRRRRRRRRVRFRC0ER0lNENCl0NHODkRVMHO0FRM#00ENRCNsRsbN0VRFRH0E#0R#NNM8s-8
-RRRRRRRRRRRRsRRCCbs#0CMRC0ERsVFlRND#NClMO0H#VRFRC0ERbHlDCClM00NHRFMF0VRE-C
-RRRRRRRRRRRRvRRq_a]BumvpR Xb	NONRoC8DCON0sNH3FMRERaCkRbs#bFCVRFRC0E
R--RRRRRRRRRRRRRavq]m_Bv upXNRbOo	NCFRL8H$R#FR0RFbsPCH8RoNRkCH8DCHMRsVF
R--RRRRRRRRRRRRRbHlDCClM00NH#FMRR0FPHCsV0$REsCHRbHlDCClM00NHRFMFvVRq_a]Bumvp3 X
R--RRRRRRRRRRRRRFaFDCR8PFCDb#CsR$lNRFOEFR#C0HFRlCbDl0CMRC0ERObN	CNoR8LF$MRH
R--RRRRRRRRRRRRRC0ER#lF0VRCVHHOCRM0lMNMCNsRPDNHNCLDRR0F0lEC3-
-
R--------------------------------------------------------------------------------
-RseC#MHFRRRR:3R46-
-R07NCRRRRRRR:cR.RDKk$gR4g-n
--R--------------------------------------------------------------------------
--
Ck#R)Wmiq3va)]_ 3qpN;DD
ObN	CNoRavq]m_Bv upX#RH
RRRRMOF#M0N0FRBbH$)ohE0FO0HC1:Rah)QtR
RRRRR:"=RB$FbsEHo0gR4gQnR 3  RDqDRosHER0#sCC#s8PC3
";
RRRR
--RRRR-a-R$RbC7HCVMHH0F
M#RRRR-R-
R0RR$RbCBumvpR XHR#
RRRRRsRRCsOF8R
RRRRRRRRRRRRRR R): R)qRp;RRRRR-RR-CR)NbDRN
s0RRRRRRRRRRRRRRRRQRv:)p q;RRRRRRRRR--QolNHsMN$NRbsR0
RRRRRCRRMs8RCsOF8
;
RRRR#0kL$RbCuQm1a Qe_q) p#RHRq) pNRsMRoCjR3j0)FR 'qp]]Qt;R

R#RRk$L0buCR)BQhQpuq_peqzH R# R)qspRNCMoRq-vau]_QFR0Ravq]Q_u;R

R0RR$RbCBumvp_ Xuqmp)#RH
RRRRRRRROsCF
s8RRRRRRRRRRRRRRRRv:qtR1umQeaQ  _)qRp;R-RR-NRvo0MHk
8CRRRRRRRRRRRRRRRRq:)tRQu)huBQqep_q pz;-RR-MRqoRDCHsMRNN8HMR#;-avq]Q_uRRH#HCDDo
NDRRRRRRRRCRM8sFCOs
8;
RRRR
--RRRR-B-RF0M#NRM07HCVMHH0F
M#RRRR-R-
RORRF0M#NRM0Ravq]A_Bq_1 4B:Rmpvu :XR=mRBv upX4'53Rj,j23j;R
RRFROMN#0MR0Rv]qa_qBA1K _:mRBv upX=R:RvBmuXp '35jj4,R3;j2
RRRRMOF#M0N0vRRq_a]B)Z mB:Rmpvu :XR=mRBv upXj'53Rj,j23j;


RRRR-R-
R-RR-PRmCFsDN88CRkCJN0DH$MRN8MRHCNJkD$H0RCFbsFN0sV#RFBsRmpvu uX_m)pq
RRRRR--5kCJN0DH$MRN8MRHCNJkD$H0RCFbsFN0sV#RFBsRmpvu NXRsbCRsCC8VCHM8R2
R-RR-R

RVRRk0MOHRFM""/=Rp5R:MRHRvBmuXp _pumqR);RR):HBMRmpvu uX_m)pqRs2RCs0kMmRAmqp hR;
RRRRR-RR-kRus#bFCR:
RRRRR-RR-RRRRRRRRCR)0Mks#)RazH RVRRpHM#RFC0RJDkNRR0F)MRN8CRs0Mks#qRwp
1 RRRRRRRR-R-RRRRRRFRR0sECICH#
RRRRRRRRR--1ObCHRNDPkNDC
#:RRRRRRRR-R-RRRRRRBRRmpvu uX_m)pq'35jjX,R2=R/RvBmuXp _pumq5)'j,3jRRY2skC0s
M#RRRRRRRR-R-RRRRRRwRRq p1RosCNDs8CR##F0VREPCRNCDkRRFVXMRN83RY
RRRRRRRRR--7NFlH
M:RRRRRRRR-R-RRRRRRpRRRRHMBumvp_ Xuqmp)MRN83RpqR)t/-=Rv]qa_
uQRRRRRRRR-R-RRRRRR)RRRRHMBumvp_ Xuqmp)MRN83R)qR)t/-=Rv]qa_
uQRRRRRRRR- -RsssFRMOF8HH0F:M#
RRRRRRRRR--RRRRRRRR FsssVRHRqp3)=tRRq-vau]_QR
RRRRRR-R-RRRRRRRRRs sFHsRV3R)qR)t=vR-q_a]uRQ
RRRRR-RR-NR)M:oC
RRRRRRRRR--RRRRRRRR""/=5)p,2#RHR0CHERCsa )zRRFsw1qp R
RRRRRR-R-R0hFC
#:RRRRRRRR-R-RRRRRRhRRF
MC
RRRRMVkOF0HM=R""RR5pH:RMmRBv upXm_up;q)R:R)RRHMBumvp_ Xuqmp)RR2skC0sAMRm mpq
h;RRRRRRRR-u-RkFsb#
C:RRRRRRRR-R-RRRRRR)RRCs0kMa#R)Rz HpVRRRH#CNJkDFR0RN)RMs8RCs0kMw#Rq p1REF0CHsI#RC
RRRRR-RR-bR1CNOHDNRPD#kC:R
RRRRRR-R-RRRRRRRRRvBmuXp _pumq5)'j,3jRRX2=mRBv upXm_up'q)5jj3,2RYR0sCk#sMRza) R
RRRRRR-R-RRRRRRRRRosCNDs8CR##F0VREPCRNCDkRRFVXMRN83RY
RRRRRRRRR--7NFlH
M:RRRRRRRR-R-RRRRRRpRRRRHMBumvp_ Xuqmp)MRN83RpqR)t/-=Rv]qa_
uQRRRRRRRR-R-RRRRRR)RRRRHMBumvp_ Xuqmp)MRN83R)qR)t/-=Rv]qa_
uQRRRRRRRR- -RsssFRMOF8HH0F:M#
RRRRRRRRR--RRRRRRRR FsssVRHRqp3)=tRRq-vau]_QR
RRRRRR-R-RRRRRRRRRs sFHsRV3R)qR)t=vR-q_a]uRQ
RRRRR-RR-NR)M:oC
RRRRRRRRR--RRRRRRRR"5="p2,)RRH#CEH0CasR)Rz FwsRq p1
RRRRRRRRR--hCF0#R:
RRRRR-RR-RRRRRRRRFRhM
C
RRRR-R-
R-RR-kRwMHO0F7MRCNODsHN0F
M#RRRR-R-
RVRRk0MOHRFMt_ auh)QBqQupq_ep5z XH:RM R)q2pRR0sCkRsMuh)QBqQupq_ep;z 
RRRRRRRRR--ubksF:#C
RRRRRRRRR--RRRRRRRR)kC0sRM#bMsHONHbDNRPDRkCFNVRMCoDRRX;XMRHR8sNH#NM
RRRRRRRRR--1ObCHRNDPkNDC
#:RRRRRRRR-R-RRRRRRhRRF
MCRRRRRRRR-7-RFHlNMR:
RRRRR-RR-RRRRRRRRRRXH)MR 
qpRRRRRRRR- -RsssFRMOF8HH0F:M#
RRRRRRRRR--RRRRRRRRhCFM
RRRRRRRRR--)oNMCR:
RRRRR-RR-RRRRRRRRvR-q_a]u<QRRat _Qu)huBQqep_q pz5RX2<v=Rq_a]uRQ
RRRRR-RR-FRh0:C#
RRRRRRRRR--RRRRRRRRhCFM
R
RRkRVMHO0FBMRvXup5RX:H)MR ;qpR:RYRRHM)p q:j=R32jRR0sCkRsMBumvp; X
RRRRRRRRR--ubksF:#C
RRRRRRRRR--RRRRRRRR)kC0sRM#BumvpR XMLklCXsRRH+RYR
RRRRRR-R-RC1bODHNRDPNk:C#
RRRRRRRRR--RRRRRRRRhCFM
RRRRRRRRR--7NFlH
M:RRRRRRRR-R-RRRRRRXRRRRHM)p q
RRRRRRRRR--RRRRRRRRYMRHRq) pR
RRRRRR-R-Rs sFOsRFHM80MHF#R:
RRRRR-RR-RRRRRRRRFRhMRC
RRRRR-RR-NR)M:oC
RRRRRRRRR--RRRRRRRRBpvuX,5XYH2R#NRl0lECNO0HN$DDRLkMF8kMCR8
RRRRR-RR-FRh0:C#
RRRRRRRRR--RRRRRRRRhCFM
R
RRkRVMHO0FuMRm)pq__amBumvp5 XZH:RMmRBv upXm_upRq)2CRs0MksRvBmuXp ;R
RRRRRR-R-RsukbCF#:R
RRRRRR-R-RRRRRRRRR0)Ck#sMRvBmuXp RDPNkFCRV
RZRRRRRRRR-1-RbHCONPDRNCDk#R:
RRRRR-RR-RRRRRRRRFRhMRC
RRRRR-RR-FR7lMNH:R
RRRRRR-R-RRRRRRRRRHZRMmRBv upXm_upRq)NRM8Z)3qt=R/Rq-vau]_QR
RRRRRR-R-Rs sFOsRFHM80MHF#R:
RRRRR-RR-RRRRRRRRsR sRFsHZVR3tq)R-=Rv]qa_
uQRRRRRRRR-)-RNCMo:R
RRRRRR-R-RRRRRRRRRpumqa)_mm_Bv upX25ZRRH#lEN0C0lNHDONDk$RMkLFM88C
RRRRRRRRR--hCF0#R:
RRRRR-RR-RRRRRRRRFRhM
C
RRRRVOkM0MHFRvBmuXp __amuqmp):5ZRRHMBumvpR X2CRs0MksRvBmuXp _pumq
);RRRRRRRR-u-RkFsb#
C:RRRRRRRR-R-RRRRRR)RRCs0kMb#RsOHMHDbNRDPNkBCRmpvu uX_m)pqRRFVZR
RRRRRR-R-RC1bODHNRDPNk:C#
RRRRRRRRR--RRRRRRRRBumvp_ Xaum_m)pq5avq]Z_B 2)mRB=Rmpvu uX_m)pq'35jjj,R3
j2RRRRRRRR-R-RRRRRRBRRmpvu aX_mm_up5q)Z=2RRvBmuXp _pumq5)'q5A1Zv3Q2R,
RRRRR-RR-RRRRRRRRRRRRRRRRRRRRRRRRRRRR1RRQ5thZv3Q2q*vau]_Qe_m .)_2VRHR)Z3 RR=j
3jRRRRRRRR-7-RFHlNMR:
RRRRR-RR-RRRRRRRRRRZHBMRmpvu RX
RRRRR-RR-sR sRFsO8FMHF0HM
#:RRRRRRRR-R-RRRRRRhRRF
MCRRRRRRRR-)-RNCMo:R
RRRRRR-R-RRRRRRRRR#sCk3D0vRqt>j=R3Rj
RRRRR-RR-RRRRRRRRvR-q_a]u<QRR#sCk3D0qR)t<v=Rq_a]uRQ
RRRRR-RR-FRh0:C#
RRRRRRRRR--RRRRRRRRhCFM
R
RRkRVMHO0F"MRq"A15RZ:HBMRmpvu uX_m)pqRs2RCs0kMmRu1QQae) _ ;qp
RRRRRRRRR--ubksF:#C
RRRRRRRRR--RRRRRRRR)kC0sRM#NFL#DCk0RDPNk5CRlMNoH80kCF2RV
RZRRRRRRRR-1-RbHCONPDRNCDk#R:
RRRRR-RR-RRRRRRRRFRhMRC
RRRRR-RR-FR7lMNH:R
RRRRRR-R-RRRRRRRRRHZRMmRBv upXm_upRq)NRM8Z)3qt=R/Rq-vau]_QR
RRRRRR-R-Rs sFOsRFHM80MHF#R:
RRRRR-RR-RRRRRRRRsR sRFsHZVR3tq)R-=Rv]qa_
uQRRRRRRRR-)-RNCMo:R
RRRRRR-R-RRRRRRRRR1qA5RZ2>j=R3Rj
RRRRR-RR-FRh0:C#
RRRRRRRRR--RRRRRRRRq5A1Z=2RRvZ3q
t
RRRRVOkM0MHFRA"q1Z"5:MRHRvBmuXp Rs2RCs0kMmRu1QQae) _ ;qp
RRRRRRRRR--ubksF:#C
RRRRRRRRR--RRRRRRRR)kC0sRM#NFL#DCk0RDPNk5CRlMNoH80kCF2RV
RZRRRRRRRR-1-RbHCONPDRNCDk#R:
RRRRR-RR-RRRRRRRRFRhMRC
RRRRR-RR-FR7lMNH:R
RRRRRR-R-RRRRRRRRRHZRMmRBv upXR
RRRRRR-R-Rs sFOsRFHM80MHF#R:
RRRRR-RR-RRRRRRRRFRhMRC
RRRRR-RR-NR)M:oC
RRRRRRRRR--RRRRRRRRq5A1ZH2R#NRl0lECNO0HN$DDRLkMF8kMCR8
RRRRR-RR-FRh0:C#
RRRRRRRRR--RRRRRRRRq5A1Z=2RR)1Ta35Z)Z *3R) +3RZQZv*32Qv
R
RRkRVMHO0FqMR)Zt5:MRHRvBmuXp _pumq2)RR0sCkRsMuh)QBqQupq_ep;z 
RRRRRRRRR--ubksF:#C
RRRRRRRRR--RRRRRRRR)kC0sRM#Nksol0CMRM5No2DCRRHMsHN8NRM#F0VREbCRsOHMHDbN
RRRRRRRRR--RRRRRRRRPkNDCVRFRRZ
RRRRR-RR-bR1CNOHDNRPD#kC:R
RRRRRR-R-RRRRRRRRRMhFCR
RRRRRR-R-Rl7FN:HM
RRRRRRRRR--RRRRRRRRZMRHRvBmuXp _pumqN)RMZ8R3tq)RR/=-avq]Q_u
RRRRRRRRR-- FsssFROM08HH#FM:R
RRRRRR-R-RRRRRRRRRs sFHsRV3RZqR)t=vR-q_a]uRQ
RRRRR-RR-NR)M:oC
RRRRRRRRR--RRRRRRRR-avq]Q_uRq<R)Zt52=R<Ravq]Q_u
RRRRRRRRR--hCF0#R:
RRRRR-RR-RRRRRRRR)Rqt25ZRZ=R3tq)
R

RVRRk0MOHRFMq5)tZH:RMmRBv upXRR2skC0suMR)BQhQpuq_peqz
 ;RRRRRRRR-u-RkFsb#
C:RRRRRRRR-R-RRRRRR)RRCs0kMN#RslokCRM05oNMDRC2HsMRNN8HMF#RVER0CsRbHHMOb
NDRRRRRRRR-R-RRRRRRPRRNCDkRRFVZR
RRRRRR-R-RC1bODHNRDPNk:C#
RRRRRRRRR--RRRRRRRRq5)tZ=2RRjj3RRHVZ 3)RR>=jR3jNRM8Zv3QRj=R3Rj
RRRRR-RR-RRRRRRRR)Rqt25ZR1=RQ5thZv3Q2q*vau]_Qe_m .)_RRHVZ 3)Rj=R3Rj
RRRRR-RR-RRRRRRRR)Rqt25ZRv=Rq_a]uHQRV3RZ)< RRjj3RRRRRRRRNRM8Zv3QRj=R3Rj
RRRRR-RR-FR7lMNH:R
RRRRRR-R-RRRRRRRRRHZRMmRBv upXR
RRRRRR-R-Rs sFOsRFHM80MHF#R:
RRRRR-RR-RRRRRRRRFRhMRC
RRRRR-RR-NR)M:oC
RRRRRRRRR--RRRRRRRR-avq]Q_uRq<R)Zt52=R<Ravq]Q_u
RRRRRRRRR--hCF0#R:
RRRRR-RR-RRRRRRRR)Rqt25ZRq=R)qBah35ZQRv,Z 3)2R

RVRRk0MOHRFM"R-"5RZ:HBMRmpvu uX_m)pqRs2RCs0kMmRBv upXm_up;q)
RRRRRRRRR--ubksF:#C
RRRRRRRRR--RRRRRRRR)kC0sRM#bMsHONHbDNRPDRkCFkVRM$NsRMlHkF#RV
RZRRRRRRRR-1-RbHCONPDRNCDk#R:
RRRRR-RR-RRRRRRRR-R""25ZRB=Rmpvu uX_m)pq'35Zv,qtRavq]Q_u2VRHRqZ3)=tRRjj3
RRRRRRRRR--7NFlH
M:RRRRRRRR-R-RRRRRRZRRRRHMBumvp_ Xuqmp)MRN83RZqR)t/-=Rv]qa_
uQRRRRRRRR- -RsssFRMOF8HH0F:M#
RRRRRRRRR--RRRRRRRR FsssVRHRqZ3)=tRRq-vau]_QR
RRRRRR-R-RM)No
C:RRRRRRRR-R-RRRRRRsRRCD#k0q3vt=R>Rjj3
RRRRRRRRR--RRRRRRRR-avq]Q_uRs<RCD#k0)3qt=R<Ravq]Q_u
RRRRRRRRR--hCF0#R:
RRRRR-RR-RRRRRRRRCR)0Mks#mRBv upXm_up'q)5vZ3qRt,Z)3qtRR-1hQt5qZ3)*t2v]qa_2uQR
HVRRRRRRRR-R-RRRRRRRRRRRRRR3RZqR)t/j=R3
j
RRRRVOkM0MHFR""-R:5ZRRHMBumvpR X2CRs0MksRvBmuXp ;R
RRRRRR-R-RsukbCF#:R
RRRRRR-R-RRRRRRRRR0)Ck#sMRNkMsl$RH#MkRRFVZR
RRRRRR-R-RC1bODHNRDPNk:C#
RRRRRRRRR--RRRRRRRRhCFM
RRRRRRRRR--7NFlH
M:RRRRRRRR-R-RRRRRRZRRRRHMBumvp
 XRRRRRRRR- -RsssFRMOF8HH0F:M#
RRRRRRRRR--RRRRRRRRhCFM
RRRRRRRRR--)oNMCR:
RRRRR-RR-RRRRRRRR-R""25ZRRH#lEN0C0lNHDONDk$RMkLFM88C
RRRRRRRRR--hCF0#R:
RRRRR-RR-RRRRRRRRCR)0Mks#GR-R$-[RsVFRRZ=GRR+[
$
RRRRVOkM0MHFRhBmKZR5:MRHRvBmuXp _pumqR)2skC0sBMRmpvu uX_m)pq;R
RRRRRR-R-RsukbCF#:R
RRRRRR-R-RRRRRRRRR0)Ck#sMRHbsMbOHNPDRNCDkRRFVObFlDRCGO[FMk0oNCVRFRRZ
RRRRR-RR-bR1CNOHDNRPD#kC:R
RRRRRR-R-RRRRRRRRRhBmK25ZRB=Rmpvu uX_m)pq'35Zv,qtRavq]Q_u2VRHRqZ3)=tRRavq]Q_u
RRRRRRRRR--7NFlH
M:RRRRRRRR-R-RRRRRRZRRRRHMBumvp_ Xuqmp)MRN83RZqR)t/-=Rv]qa_
uQRRRRRRRR- -RsssFRMOF8HH0F:M#
RRRRRRRRR--RRRRRRRR FsssVRHRqZ3)=tRRq-vau]_QR
RRRRRR-R-RM)No
C:RRRRRRRR-R-RRRRRRsRRCD#k0q3vt=R>Rjj3
RRRRRRRRR--RRRRRRRR-avq]Q_uRs<RCD#k0)3qt=R<Ravq]Q_u
RRRRRRRRR--hCF0#R:
RRRRR-RR-RRRRRRRRCR)0Mks#mRBv upXm_up'q)5vZ3qRt,-qZ3)Rt2HZVR3tq)RR/=v]qa_
uQ
RRRRMVkOF0HMmRBh5KRZH:RMmRBv upXs2RCs0kMmRBv upXR;
RRRRR-RR-kRus#bFCR:
RRRRR-RR-RRRRRRRRCR)0Mks#FROlCbDGFROMo[kNR0CFZVR
RRRRRRRRR--1ObCHRNDPkNDC
#:RRRRRRRR-R-RRRRRRhRRF
MCRRRRRRRR-7-RFHlNMR:
RRRRR-RR-RRRRRRRRRRZHBMRmpvu RX
RRRRR-RR-sR sRFsO8FMHF0HM
#:RRRRRRRR-R-RRRRRRhRRF
MCRRRRRRRR-)-RNCMo:R
RRRRRR-R-RRRRRRRRRhBmK25ZRRH#lEN0C0lNHDONDk$RMkLFM88C
RRRRRRRRR--hCF0#R:
RRRRR-RR-RRRRRRRRCR)0Mks#RRG-R[$VRFsZG=RR[+R$R

RVRRk0MOHRFM1aT)5RZ:HBMRmpvu uX_m)pqRs2RCs0kMmRBv upXm_up;q)
RRRRRRRRR--ubksF:#C
RRRRRRRRR--RRRRRRRR)kC0sRM##NJkssCRFRF0FZVRR0IHEFRb#HH0PsCRCRNDb0Ns
RRRRRRRRR--RRRRRRRRFRs,H0VREsCRCRNDb0NsRRH#xFCs,ER0CMRFCHRI0MERFCMMoHN0PRC
RRRRR-RR-RRRRRRRRlRHNMoHNRs$b0Ns
RRRRRRRRR--1ObCHRNDPkNDC
#:RRRRRRRR-R-RRRRRR1RRT5)aZ=2RRvBmuXp _pumq5)'j,3jRjj32VRHRvZ3q=tRRjj3
RRRRRRRRR--7NFlH
M:RRRRRRRR-R-RRRRRRZRRRRHMBumvp_ Xuqmp)MRN83RZqR)t/-=Rv]qa_
uQRRRRRRRR- -RsssFRMOF8HH0F:M#
RRRRRRRRR--RRRRRRRR FsssVRHRqZ3)=tRRq-vau]_QR
RRRRRR-R-RM)No
C:RRRRRRRR-R-RRRRRRsRRCD#k0q3vt=R>Rjj3
RRRRRRRRR--RRRRRRRR-avq]Q_uRs<RCD#k0)3qt=R<Ravq]Q_u
RRRRRRRRR--hCF0#R:
RRRRR-RR-RRRRRRRRFRhM
C
RRRRVOkM0MHFR)1Ta:5ZRRHMBumvpR X2CRs0MksRvBmuXp ;R
RRRRRR-R-RsukbCF#:R
RRRRRR-R-RRRRRRRRR0)Ck#sMRk#JNRsCs0FFRRFVZHRI0bERF0#HHRPCsDCNRsbN0R
RRRRRR-R-RRRRRRRRR,FsRRHV0RECsDCNRsbN0#RHRsxCF0,REFCRMICRHR0EMMFMC0oNH
PCRRRRRRRR-R-RRRRRRHRRlHNoM$NsRsbN0R
RRRRRR-R-RC1bODHNRDPNk:C#
RRRRRRRRR--RRRRRRRR1aT)5avq]Z_B 2)mRv=Rq_a]B)Z mR
RRRRRR-R-Rl7FN:HM
RRRRRRRRR--RRRRRRRRZMRHRvBmuXp 
RRRRRRRRR-- FsssFROM08HH#FM:R
RRRRRR-R-RRRRRRRRRMhFCR
RRRRRR-R-RM)No
C:RRRRRRRR-R-RRRRRR1RRT5)aZH2R#NRl0lECNO0HN$DDRLkMF8kMCR8
RRRRR-RR-FRh0:C#
RRRRRRRRR--RRRRRRRRhCFM
R
RRkRVMHO0F MRXZu5:MRHRvBmuXp _pumq2)RR0sCkRsMBumvp_ Xuqmp)R;
RRRRR-RR-kRus#bFCR:
RRRRR-RR-RRRRRRRRCR)0Mks#sRbHHMObRNDPkNDCVRFRbCGFMMC0DHNRRFVZR
RRRRRR-R-RC1bODHNRDPNk:C#
RRRRRRRRR--RRRRRRRR 5XuZ=2RRvBmuXp _pumq5)'4,3jRjj32VRHRvZ3q=tRjR3jN
M8RRRRRRRR-R-RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR3RZqR)t=3RjjR
RRRRRR-R-RRRRRRRRRu X5RZ2=mRBv upXm_up'q)5j43,qRvau]_QH2RV3RZvRqt=qRvau]_QMRN8R
RRRRRR-R-RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRq5A1Z)3qt=2RRavq]Q_u_ me)
_.RRRRRRRR-R-RRRRRR RRXZu52RR=Bumvp_ Xuqmp)4'53Rj,v]qa__uQm)e _R.2HRV
RRRRR-RR-RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRvZ3q=tRRavq]Q_u_ me)R_.N
M8RRRRRRRR-R-RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR3RZqR)t=qRvau]_Qe_m .)_
RRRRRRRRR--RRRRRRRR 5XuZ=2RRvBmuXp _pumq5)'4,3jRq-vau]_Qe_m .)_2VRH
RRRRRRRRR--RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRZRR3tvqRv=Rq_a]umQ_e_ ).MRN8R
RRRRRR-R-RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRZ)3qtRR=-avq]Q_u_ me)
_.RRRRRRRR-7-RFHlNMR:
RRRRR-RR-RRRRRRRRRRZHBMRmpvu uX_m)pqR8NMRqZ3)/tR=vR-q_a]uRQ
RRRRR-RR-sR sRFsO8FMHF0HM
#:RRRRRRRR-R-RRRRRR RRsssFRRHVZ)3qtRR=-avq]Q_u
RRRRRRRRR--)oNMCR:
RRRRR-RR-RRRRRRRRCRs#0kD3tvqRR>=j
3jRRRRRRRR-R-RRRRRR-RRv]qa_RuQ<CRs#0kD3tq)RR<=v]qa_
uQRRRRRRRR-h-RF#0C:R
RRRRRR-R-RRRRRRRRRMhFCR

RVRRk0MOHRFM 5XuZH:RMmRBv upXRR2skC0sBMRmpvu 
X;RRRRRRRR-u-RkFsb#
C:RRRRRRRR-R-RRRRRR)RRCs0kMC#RGMbFCHM0NFDRV
RZRRRRRRRR-1-RbHCONPDRNCDk#R:
RRRRR-RR-RRRRRRRRXR uq5vaB]_Zm )2RR=v]qa_qBA14 _
RRRRRRRRR--RRRRRRRR 5XuZ=2RRq-vaB]_A q1_H4RV3RZ)= RRjj3R8NMR1qA5QZ3v=2RRavq]Q_u
RRRRRRRRR--RRRRRRRR 5XuZ=2RRt1Qh35ZQ*v2v]qa_qBA1K _RRHVZ 3)Rj=R3NjRMR8
RRRRR-RR-RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRqRRAZ1532QvRR=Rv]qa__uQm)e _R.
RRRRR-RR-FR7lMNH:R
RRRRRR-R-RRRRRRRRRHZRMmRBv upXR
RRRRRR-R-Rs sFOsRFHM80MHF#R:
RRRRR-RR-RRRRRRRRFRhMRC
RRRRR-RR-NR)M:oC
RRRRRRRRR--RRRRRRRR 5XuZH2R#NRl0lECNO0HN$DDRLkMF8kMCR8
RRRRR-RR-FRh0:C#
RRRRRRRRR--RRRRRRRRhCFM



RRRRVOkM0MHFRtpm.:5ZRRHMBumvpR X2CRs0MksRvBmuXp ;R
RRRRRR-R-RsukbCF#:R
RRRRRR-R-RRRRRRRRR0)Ck#sMRoDFN0sHELlRNR#C.VRFRRZ
RRRRR-RR-bR1CNOHDNRPD#kC:R
RRRRRR-R-RRRRRRRRRtpm.q5vaB]_A q1_R42=qRvaB]_Zm )
RRRRRRRRR--RRRRRRRRp.mt5RZ2=qRvaB]_A q1_H4RVRRZ=mRBv upX.'53Rj,j23j
RRRRRRRRR--7NFlH
M:RRRRRRRR-R-RRRRRRZRRRRHMBumvpR XNRM8q5A1Z/2R=3RjjR
RRRRRR-R-Rs sFOsRFHM80MHF#R:
RRRRR-RR-RRRRRRRRsR sRFsHqVRAZ152RR=j
3jRRRRRRRR-)-RNCMo:R
RRRRRR-R-RRRRRRRRRtpm.25ZRRH#lEN0C0lNHDONDk$RMkLFM88C
RRRRRRRRR--hCF0#R:
RRRRR-RR-RRRRRRRRFRhM
C
RRRRVOkM0MHFRtpm5RZ:HBMRmpvu 2XRR0sCkRsMBumvp; X
RRRRRRRRR--ubksF:#C
RRRRRRRRR--RRRRRRRR)kC0sRM#MkN0sRNDDNFosEH0lVRFRRZ
RRRRR-RR-bR1CNOHDNRPD#kC:R
RRRRRR-R-RRRRRRRRRtpm5avq]A_Bq_1 4=2RRavq]Z_B 
)mRRRRRRRR-R-RRRRRRpRRm-t5v]qa_qBA14 _2RR=Bumvp' X5jj3,qRvau]_QR2
RRRRR-RR-RRRRRRRRmRptq5vaB]_A q1_RK2=mRBv upXj'53Rj,v]qa__uQm)e _
.2RRRRRRRR-R-RRRRRRpRRm-t5v]qa_qBA1K _2RR=Bumvp' X5jj3,vR-q_a]umQ_e_ ).R2
RRRRR-RR-RRRRRRRRmRpt25ZRv=Rq_a]B1Aq R_4HZVRRB=Rmpvu 5X'v]qa_R ,j23j
RRRRRRRRR--7NFlH
M:RRRRRRRR-R-RRRRRRZRRRRHMBumvpR XNRM8q5A1Z/2R=3RjjR
RRRRRR-R-Rs sFOsRFHM80MHF#R:
RRRRR-RR-RRRRRRRRsR sRFsHqVRAZ152RR=j
3jRRRRRRRR-)-RNCMo:R
RRRRRR-R-RRRRRRRRRtpm5RZ2Hl#RNC0ElHN0ODND$MRkLMFk8
C8RRRRRRRR-h-RF#0C:R
RRRRRR-R-RRRRRRRRRMhFCR

RVRRk0MOHRFMp4mtj:5ZRRHMBumvpR X2CRs0MksRvBmuXp ;R
RRRRRR-R-RsukbCF#:R
RRRRRR-R-RRRRRRRRR0)Ck#sMRoDFN0sHELlRNR#C4FjRV
RZRRRRRRRR-1-RbHCONPDRNCDk#R:
RRRRR-RR-RRRRRRRRmRpt54jv]qa_qBA14 _2RR=v]qa_ BZ)Rm
RRRRR-RR-RRRRRRRRmRpt54jZ=2RRavq]A_Bq_1 4VRHR=ZRRvBmuXp 'j543Rj,j23j
RRRRRRRRR--7NFlH
M:RRRRRRRR-R-RRRRRRZRRRRHMBumvpR XNRM8q5A1Z/2R=3RjjR
RRRRRR-R-Rs sFOsRFHM80MHF#R:
RRRRR-RR-RRRRRRRRsR sRFsHqVRAZ152RR=j
3jRRRRRRRR-)-RNCMo:R
RRRRRR-R-RRRRRRRRRtpm4Zj52#RHR0lNENCl0NHODRD$kFMLkCM88R
RRRRRR-R-R0hFC
#:RRRRRRRR-R-RRRRRRhRRF
MC
RRRRMVkOF0HMmRptZ.5:MRHRvBmuXp _pumq2)RR0sCkRsMBumvp_ Xuqmp)R;
RRRRR-RR-kRus#bFCR:
RRRRR-RR-RRRRRRRRCR)0Mks#sRbHHMObRNDPkNDCVRFRoDFN0sHELlRNR#C.VRFRRZ
RRRRR-RR-bR1CNOHDNRPD#kC:R
RRRRRR-R-RRRRRRRRRtpm.25ZRB=Rmpvu uX_m)pq'35jjj,R3Rj2HZVR3tvqR4=R3NjRMR8
RRRRR-RR-RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRZRR3tq)Rj=R3Rj
RRRRR-RR-RRRRRRRRmRptZ.52RR=Bumvp_ Xuqmp)4'53Rj,j23jRRHVZq3vtRR=.R3jN
M8RRRRRRRR-R-RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRZRR3tq)Rj=R3Rj
RRRRR-RR-FR7lMNH:R
RRRRRR-R-RRRRRRRRRHZRMmRBv upXm_upRq)NRM8Z)3qt=R/Rq-vau]_QR
RRRRRR-R-RRRRRRRRRvZ3q/tR=3RjjR
RRRRRR-R-Rs sFOsRFHM80MHF#R:
RRRRR-RR-RRRRRRRRsR sRFsHZVR3tq)R-=Rv]qa_
uQRRRRRRRR-R-RRRRRR RRsssFRRHVZq3vtRR=j
3jRRRRRRRR-)-RNCMo:R
RRRRRR-R-RRRRRRRRR#sCk3D0vRqt>j=R3Rj
RRRRR-RR-RRRRRRRRvR-q_a]u<QRR#sCk3D0qR)t<v=Rq_a]uRQ
RRRRR-RR-FRh0:C#
RRRRRRRRR--RRRRRhRRF
MC
RRRRMVkOF0HMmRpt:5ZRRHMBumvp_ Xuqmp)RR2skC0sBMRmpvu uX_m)pq;R
RRRRRR-R-RsukbCF#:R
RRRRRR-R-RRRRRRRRR0)Ck#sMRHbsMbOHNPDRNCDkRRFVMkN0sRNDDNFosEH0lVRFRRZ
RRRRR-RR-bR1CNOHDNRPD#kC:R
RRRRRR-R-RRRRRRRRRtpm5RZ2=mRBv upXm_up'q)5jj3,3RjjH2RV3RZvRqt=3R4jMRN8R
RRRRRR-R-RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRqZ3)=tRRjj3
RRRRRRRRR--RRRRRRRRp5mtZ=2RRvBmuXp _pumq5)'v]qa_,uQRavq]Q_u_ me)2_.R
HVRRRRRRRR-R-RRRRRRRRRRRRRRRRRRRRRRRRRRRRRZq3vtRR=4R3jNRM8Z)3qtRR=v]qa_
uQRRRRRRRR-R-RRRRRRpRRmZt52RR=Bumvp_ Xuqmp)v'5q_a]umQ_e_ ).v,Rq_a]umQ_e_ ).H2RVR
RRRRRR-R-RRRRRRRRRRRRRRRRRRRRRRRRRRRRR3RZvRqt=3R4jMRN8ZRR3tq)Rv=Rq_a]umQ_e_ ).R
RRRRRR-R-RRRRRRRRRtpm5RZ2=mRBv upXm_up'q)5avq]Q_u_ me),_.Rq-vau]_Qe_m .)_2VRH
RRRRRRRRR--RRRRRRRRRRRRRRRRRRRRRRRRRRRRRvZ3q=tRRj43R8NMR3RZqR)t=vR-q_a]umQ_e_ ).R
RRRRRR-R-RRRRRRRRRtpm5RZ2=mRBv upXm_up'q)5j43,3RjjH2RV3RZvRqt=qRva ]_R8NM
RRRRRRRRR--RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRZ)3qtRR=j
3jRRRRRRRR-7-RFHlNMR:
RRRRR-RR-RRRRRRRRRRZHBMRmpvu uX_m)pqR8NMRqZ3)/tR=vR-q_a]uRQ
RRRRR-RR-RRRRRRRR3RZvRqt/j=R3Rj
RRRRR-RR-sR sRFsO8FMHF0HM
#:RRRRRRRR-R-RRRRRR RRsssFRRHVZ)3qtRR=-avq]Q_u
RRRRRRRRR--RRRRRRRR FsssVRHRvZ3q=tRRjj3
RRRRRRRRR--)oNMCR:
RRRRR-RR-RRRRRRRRCRs#0kD3tvqRR>=j
3jRRRRRRRR-R-RRRRRR-RRv]qa_RuQ<CRs#0kD3tq)RR<=v]qa_
uQRRRRRRRR-h-RF#0C:R
RRRRRR-R-RRRRRRRRRMhFCR

RVRRk0MOHRFMp4mtj:5ZRRHMBumvp_ Xuqmp)RR2skC0sBMRmpvu uX_m)pq;R
RRRRRR-R-RsukbCF#:R
RRRRRR-R-RRRRRRRRR0)Ck#sMRHbsMbOHNPDRNCDkRRFVDNFosEH0lNRL#4CRjVRFRRZ
RRRRR-RR-bR1CNOHDNRPD#kC:R
RRRRRR-R-RRRRRRRRRtpm4Zj52RR=Bumvp_ Xuqmp)j'53Rj,j23jRRHVZq3vtRR=4R3jN
M8RRRRRRRR-R-RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRqZ3)=tRRjj3
RRRRRRRRR--RRRRRRRRp4mtj25ZRB=Rmpvu uX_m)pq'354jj,R3Rj2HZVR3tvqR4=RjR3jN
M8RRRRRRRR-R-RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRqZ3)=tRRjj3
RRRRRRRRR--7NFlH
M:RRRRRRRR-R-RRRRRRZRRRRHMBumvp_ Xuqmp)MRN83RZqR)t/-=Rv]qa_
uQRRRRRRRR-R-RRRRRRZRR3tvqRR/=j
3jRRRRRRRR- -RsssFRMOF8HH0F:M#
RRRRRRRRR--RRRRRRRR FsssVRHRqZ3)=tRRq-vau]_QR
RRRRRR-R-RRRRRRRRRs sFHsRV3RZvRqt=3RjjR
RRRRRR-R-RM)No
C:RRRRRRRR-R-RRRRRRsRRCD#k0q3vt=R>Rjj3
RRRRRRRRR--RRRRRRRR-avq]Q_uRs<RCD#k0)3qt=R<Ravq]Q_u
RRRRRRRRR--hCF0#R:
RRRRR-RR-RRRRRRRRFRhM
C
RRRRVOkM0MHFRtpm5RZ:HBMRmpvu RX;A q1:MRHRq) ps2RCs0kMmRBv upXR;
RRRRR-RR-kRus#bFCR:
RRRRR-RR-RRRRRRRRCR)0Mks#FRDoHNs0RElLCN#R1Aq VRFRRZ
RRRRR-RR-bR1CNOHDNRPD#kC:R
RRRRRR-R-RRRRRRRRRtpm5avq]A_Bq_1 4A,Rq21 Rv=Rq_a]B)Z mR
RRRRRR-R-RRRRRRRRRtpm5AZ,q21 Rv=Rq_a]B1Aq R_4HZVRRB=Rmpvu 5X'A q1,3RjjR2
RRRRR-RR-FR7lMNH:R
RRRRRR-R-RRRRRRRRRHZRMmRBv upXMRN8ARq125ZRR/=j
3jRRRRRRRR-R-RRRRRRARRqR1 >3RjjR
RRRRRR-R-RRRRRRRRR1Aq =R/Rj43
RRRRRRRRR-- FsssFROM08HH#FM:R
RRRRRR-R-RRRRRRRRRs sFHsRVARq125ZRj=R3Rj
RRRRR-RR-RRRRRRRRsR sRFsHAVRqR1 <j=R3Rj
RRRRR-RR-RRRRRRRRsR sRFsHAVRqR1 =3R4jR
RRRRRR-R-RM)No
C:RRRRRRRR-R-RRRRRRpRRmZt5,1Aq H2R#NRl0lECNO0HN$DDRLkMF8kMCR8
RRRRR-RR-FRh0:C#
RRRRRRRRR--RRRRRRRRhCFM
R
RRkRVMHO0FpMRmZt5:MRHRvBmuXp _pumqR);A q1:MRHRq) pRR2skC0sBMRmpvu uX_m)pq;R
RRRRRR-R-RsukbCF#:R
RRRRRR-R-RRRRRRRRR0)Ck#sMRHbsMbOHNPDRNCDkRRFVDNFosEH0lNRL#ACRqR1 FZVR
RRRRRRRRR--1ObCHRNDPkNDC
#:RRRRRRRR-R-RRRRRRpRRmZt5,qRA1R 2=mRBv upXm_up'q)5jj3,3RjjH2RV3RZvRqt=3R4jMRN8R
RRRRRR-R-RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRZ)3qtRR=j
3jRRRRRRRR-R-RRRRRRpRRmZt5,qRA1R 2=mRBv upXm_up'q)5j43,3RjjH2RV3RZvRqt=qRA1N RMR8
RRRRR-RR-RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRqZ3)=tRRjj3
RRRRRRRRR--7NFlH
M:RRRRRRRR-R-RRRRRRZRRRRHMBumvp_ Xuqmp)MRN83RZqR)t/-=Rv]qa_
uQRRRRRRRR-R-RRRRRRZRR3tvqRR/=j
3jRRRRRRRR-R-RRRRRRARRqR1 >3RjjR
RRRRRR-R-RRRRRRRRR1Aq =R/Rj43
RRRRRRRRR-- FsssFROM08HH#FM:R
RRRRRR-R-RRRRRRRRRs sFHsRV3RZqR)t=vR-q_a]uRQ
RRRRR-RR-RRRRRRRRsR sRFsHZVR3tvqRj=R3Rj
RRRRR-RR-RRRRRRRRsR sRFsHAVRqR1 <j=R3Rj
RRRRR-RR-RRRRRRRRsR sRFsHAVRqR1 =3R4jR
RRRRRR-R-RM)No
C:RRRRRRRR-R-RRRRRRsRRCD#k0q3vt=R>Rjj3
RRRRRRRRR--RRRRRRRR-avq]Q_uRs<RCD#k0)3qt=R<Ravq]Q_u
RRRRRRRRR--hCF0#R:
RRRRR-RR-RRRRRRRRFRhM
C
RRRRVOkM0MHFRh1QRR5Z:MRHRvBmuXp _pumq2)RR0sCkRsMBumvp_ Xuqmp)R;
RRRRR-RR-kRus#bFCR:
RRRRR-RR-RRRRRRRRCR)0Mks#sRbHHMObRNDPkNDCVRFRM#HCVRFRRZ
RRRRR-RR-bR1CNOHDNRPD#kC:R
RRRRRR-R-RRRRRRRRRh1Q5RZ2=mRBv upXm_up'q)5jj3,3RjjH2RV3RZvRqt=3RjjMRN8R
RRRRRR-R-RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRZ)3qtRR=j
3jRRRRRRRR-R-RRRRRR1RRQZh52RR=Bumvp_ Xuqmp)j'53Rj,j23jRRHVZq3vtRR=v]qa_RuQN
M8RRRRRRRR-R-RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR3RZqR)t=3RjjR
RRRRRR-R-Rl7FN:HM
RRRRRRRRR--RRRRRRRRZMRHRvBmuXp _pumqN)RMZ8R3tq)RR/=-avq]Q_u
RRRRRRRRR-- FsssFROM08HH#FM:R
RRRRRR-R-RRRRRRRRRs sFHsRV3RZqR)t=vR-q_a]uRQ
RRRRR-RR-NR)M:oC
RRRRRRRRR--RRRRRRRRskC#Dv03q>tR=3RjjR
RRRRRR-R-RRRRRRRRRq-vau]_QRR<skC#Dq03)<tR=qRvau]_QR
RRRRRR-R-R0hFC
#:RRRRRRRR-R-RRRRRRhRRF
MC
RRRRMVkOF0HMQR1hZR5RH:RMmRBv upXRR2skC0sBMRmpvu 
X;RRRRRRRR-u-RkFsb#
C:RRRRRRRR-R-RRRRRR)RRCs0kM##RHRMCFZVR
RRRRRRRRR--1ObCHRNDPkNDC
#:RRRRRRRR-R-RRRRRR1RRQvh5q_a]B)Z m=2RRavq]Z_B 
)mRRRRRRRR-R-RRRRRR1RRQZh52RR=v]qa_ BZ)HmRVRRZ=mRBv upXv'5q_a]uRQ,j23j
RRRRRRRRR--7NFlH
M:RRRRRRRR-R-RRRRRRZRRRRHMBumvp
 XRRRRRRRR- -RsssFRMOF8HH0F:M#
RRRRRRRRR--RRRRRRRRhCFM
RRRRRRRRR--)oNMCR:
RRRRR-RR-RRRRRRRRARq1Q51h25Z2=R<R)1TaQ51h35Z)* 215QhZ 3)2
R+RRRRRRRR-R-RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR1RRQ5h]Zv3Q2Q*1hZ]532Qv2R
RRRRRR-R-R0hFC
#:RRRRRRRR-R-RRRRRRhRRF
MC
RRRRMVkOF0HMBRRm51RZRR:HBMRmpvu 2XRR0sCkRsMBumvp; X
RRRRRRRRR--ubksF:#C
RRRRRRRRR--RRRRRRRR)kC0sRM#OHF#MFCRV
RZRRRRRRRR-1-RbHCONPDRNCDk#R:
RRRRR-RR-RRRRRRRRmRB125ZRv=Rq_a]B)Z mVRHR=ZRRvBmuXp 'q5vau]_Qe_m .)_,3RjjR2
RRRRR-RR-RRRRRRRRmRB125ZRv=Rq_a]B)Z mVRHR=ZRRvBmuXp 'v5-q_a]umQ_e_ ).j,R3
j2RRRRRRRR-7-RFHlNMR:
RRRRR-RR-RRRRRRRRRRZHBMRmpvu RX
RRRRR-RR-sR sRFsO8FMHF0HM
#:RRRRRRRR-R-RRRRRRhRRF
MCRRRRRRRR-)-RNCMo:R
RRRRRR-R-RRRRRRRRR1qA51Bm52Z2RR<=1aT)51Bm5)Z3 B2*mZ1532) RR+
RRRRR-RR-RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRQR1hZ]532Qv*h1Q]35ZQ2v2
RRRRRRRRR--hCF0#R:
RRRRR-RR-RRRRRRRRFRhM
C

RRRRMVkOF0HMBRRm51RZRR:HBMRmpvu uX_m)pqRs2RCs0kMmRBv upXm_up;q)
RRRRRRRRR--ubksF:#C
RRRRRRRRR--RRRRRRRR)kC0sRM#bMsHONHbDNRPDRkCFOVRFM#HCVRFRRZ
RRRRR-RR-bR1CNOHDNRPD#kC:R
RRRRRR-R-RRRRRRRRR1Bm5RZ2=mRBv upXm_up'q)5jj3,3RjjH2RV3RZvRqt=qRvau]_Qe_m .)_
RRRRRRRRR--RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRMRN83RZqR)t=3RjjR
RRRRRR-R-RRRRRRRRR1Bm5RZ2=mRBv upXm_up'q)5jj3,3RjjH2RV3RZvRqt=qRvau]_Qe_m .)_
RRRRRRRRR--RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRMRN83RZqR)t=qRvau]_QR
RRRRRR-R-Rl7FN:HM
RRRRRRRRR--RRRRRRRRZMRHRvBmuXp _pumqN)RMZ8R3tq)RR/=-avq]Q_u
RRRRRRRRR-- FsssFROM08HH#FM:R
RRRRRR-R-RRRRRRRRRs sFHsRV3RZqR)t=vR-q_a]uRQ
RRRRR-RR-NR)M:oC
RRRRRRRRR--RRRRRRRRskC#Dv03q>tR=3RjjR
RRRRRR-R-RRRRRRRRRq-vau]_QRR<skC#Dq03)<tR=qRvau]_QR
RRRRRR-R-R0hFC
#:RRRRRRRR-R-RRRRRRhRRF
MC
RRRRMVkOF0HMQR1h5]RZRR:HBMRmpvu 2XRR0sCkRsMBumvp; X
RRRRRRRRR--ubksF:#C
RRRRRRRRR--RRRRRRRR)kC0sRM#EC$bsDLFH#ORHRMCFZVR
RRRRRRRRR--1ObCHRNDPkNDC
#:RRRRRRRR-R-RRRRRR1RRQ5h]v]qa_ BZ)Rm2=qRvaB]_Zm )
RRRRRRRRR--RRRRRRRR1]Qh5RZ2=qRvaB]_Zm )RRHVZ 3)Rj=R3NjRMZ8R3RQv=qRvau]_QR
RRRRRR-R-RRRRRRRRRh1Q]25ZRv=Rq_a]B1Aq R_KHZVR3R) =3RjjMRN8R
RRRRRR-R-RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRZRR3RQv=qRvau]_Qe_m .)_
RRRRRRRRR--RRRRRRRR1]Qh5RZ2=vR-q_a]B1Aq R_KHZVR3R) =3RjjMRN8R
RRRRRR-R-RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRZRR3RQv=vR-q_a]umQ_e_ ).R
RRRRRR-R-Rl7FN:HM
RRRRRRRRR--RRRRRRRRZMRHRvBmuXp 
RRRRRRRRR-- FsssFROM08HH#FM:R
RRRRRR-R-RRRRRRRRRMhFCR
RRRRRR-R-RM)No
C:RRRRRRRR-R-RRRRRRqRRA115Q5h]ZR22<1=RT5)a1]Qh5)Z3 12*Q5h]Z 3)2
R+RRRRRRRR-R-RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR1RRQZh532Qv*h1Q5QZ3v
22RRRRRRRR-h-RF#0C:R
RRRRRR-R-RRRRRRRRRMhFCR

RVRRk0MOHRFM1]QhRR5Z:MRHRvBmuXp _pumq2)RR0sCkRsMBumvp_ Xuqmp)R;
RRRRR-RR-kRus#bFCR:
RRRRR-RR-RRRRRRRRCR)0Mks#sRbHHMObRNDPkNDCVRFRbE$CFsLDRHO#CHMRRFVZR
RRRRRR-R-RC1bODHNRDPNk:C#
RRRRRRRRR--RRRRRRRR1]Qh5RZ2=mRBv upXm_up'q)5jj3,3RjjH2RV3RZvRqt=3RjjMRN8R
RRRRRR-R-RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRZ)3qtRR=j
3jRRRRRRRR-R-RRRRRR1RRQ5h]Z=2RRvBmuXp _pumq5)'j,3jRjj32VRHRvZ3q=tRRavq]Q_uR8NM
RRRRRRRRR--RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRZRR3tq)Rv=Rq_a]umQ_e_ ).R
RRRRRR-R-RRRRRRRRRh1Q]25ZRB=Rmpvu uX_m)pq'354jv,Rq_a]umQ_e_ ).H2RV3RZvRqt=R
RRRRRR-R-RRRRRRRRRRRRRRRRRRRRRRRRRavq]Q_u_ me)R_.NRM8Z)3qtRR=v]qa__uQm)e _R.
RRRRR-RR-RRRRRRRRQR1hZ]52RR=Bumvp_ Xuqmp)4'53Rj,-avq]Q_u_ me)2_.RRHVZq3vt
R=RRRRRRRR-R-RRRRRRRRRRRRRRRRRRRRRRvRRq_a]umQ_e_ ).MRN83RZqR)t=vR-q_a]umQ_e_ ).R
RRRRRR-R-Rl7FN:HM
RRRRRRRRR--RRRRRRRRZMRHRvBmuXp _pumqN)RMZ8R3tq)RR/=-avq]Q_u
RRRRRRRRR-- FsssFROM08HH#FM:R
RRRRRR-R-RRRRRRRRRs sFHsRV3RZqR)t=vR-q_a]uRQ
RRRRR-RR-NR)M:oC
RRRRRRRRR--RRRRRRRRskC#Dv03q>tR=3RjjR
RRRRRR-R-RRRRRRRRRq-vau]_QRR<skC#Dq03)<tR=qRvau]_QR
RRRRRR-R-R0hFC
#:RRRRRRRR-R-RRRRRRhRRF
MC
RRRRMVkOF0HMmRB15]RZRR:HBMRmpvu 2XRR0sCkRsMBumvp; X
RRRRRRRRR--ubksF:#C
RRRRRRRRR--RRRRRRRR)kC0sRM#EC$bsDLFHOORFM#HCVRFRRZ
RRRRR-RR-bR1CNOHDNRPD#kC:R
RRRRRR-R-RRRRRRRRR1Bm]q5vaB]_Zm )2RR=v]qa_qBA14 _
RRRRRRRRR--RRRRRRRRB]m15RZ2=vR-q_a]B1Aq R_4HZVR3R) =3RjjMRN83RZQ=vRRavq]Q_u
RRRRRRRRR--RRRRRRRRB]m15RZ2=qRvaB]_Zm )RRHVZ 3)Rj=R3NjRMZ8R3RQv=qRvau]_Qe_m .)_
RRRRRRRRR--RRRRRRRRB]m15RZ2=qRvaB]_Zm )RRHVZ 3)Rj=R3NjRMZ8R3RQv=vR-q_a]umQ_e_ ).R
RRRRRR-R-Rl7FN:HM
RRRRRRRRR--RRRRRRRRZMRHRvBmuXp 
RRRRRRRRR-- FsssFROM08HH#FM:R
RRRRRR-R-RRRRRRRRRMhFCR
RRRRRR-R-RM)No
C:RRRRRRRR-R-RRRRRRqRRAB15m51]ZR22<1=RT5)a1]Qh5)Z3 12*Q5h]Z 3)2
R+RRRRRRRR-R-RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRBRRmZ1532Qv*1Bm5QZ3v
22RRRRRRRR-h-RF#0C:R
RRRRRR-R-RRRRRRRRRMhFC


RRRRVOkM0MHFR1Bm]ZR5RH:RMmRBv upXm_upRq)2CRs0MksRvBmuXp _pumq
);RRRRRRRR-u-RkFsb#
C:RRRRRRRR-R-RRRRRR)RRCs0kMb#RsOHMHDbNRDPNkFCRV$REbLCsFODHR#OFHRMCFZVR
RRRRRRRRR--1ObCHRNDPkNDC
#:RRRRRRRR-R-RRRRRRBRRm51]Z=2RRvBmuXp _pumq5)'4,3jRjj32VRHRvZ3q=tRRjj3R8NM
RRRRRRRRR--RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRZRR3tq)Rj=R3Rj
RRRRR-RR-RRRRRRRRmRB1Z]52RR=Bumvp_ Xuqmp)4'53Rj,v]qa_2uQRRHVZq3vtRR=v]qa_RuQN
M8RRRRRRRR-R-RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR3RZqR)t=qRvau]_Qe_m .)_
RRRRRRRRR--RRRRRRRRB]m15RZ2=mRBv upXm_up'q)5jj3,3RjjH2RV3RZvRqt=R
RRRRRR-R-RRRRRRRRRRRRRRRRRRRRRRRRv]qa__uQm)e _N.RMZ8R3tq)Rv=Rq_a]umQ_e_ ).R
RRRRRR-R-RRRRRRRRR1Bm]25ZRB=Rmpvu uX_m)pq'35jjj,R3Rj2HZVR3tvqRR=
RRRRR-RR-RRRRRRRRRRRRRRRRRRRRRRRRavq]Q_u_ me)R_.NRM8Z)3qtRR=-avq]Q_u_ me)
_.RRRRRRRR-7-RFHlNMR:
RRRRR-RR-RRRRRRRRRRZHBMRmpvu uX_m)pqR8NMRqZ3)/tR=vR-q_a]uRQ
RRRRR-RR-sR sRFsO8FMHF0HM
#:RRRRRRRR-R-RRRRRR RRsssFRRHVZ)3qtRR=-avq]Q_u
RRRRRRRRR--)oNMCR:
RRRRR-RR-RRRRRRRRCRs#0kD3tvqRR>=j
3jRRRRRRRR-R-RRRRRR-RRv]qa_RuQ<CRs#0kD3tq)RR<=v]qa_
uQRRRRRRRR-h-RF#0C:R
RRRRRR-R-RRRRRRRRRMhFCR

R-RR-R
RR-R-RHqs0CEl0RHOmsbCNs0F#R
RR-R-
R
RRkRVMHO0F"MR+5"RRRp:HBMRmpvu RX;RR):HBMRmpvu 2XRR0sCkRsMBumvp; X
RRRRRRRRR--ubksF:#C
RRRRRRRRR--RRRRRRRR)kC0sRM#N0sHE0lCHNOR808HHRFMFpVRR8NMRR)
RRRRR-RR-bR1CNOHDNRPD#kC:R
RRRRRR-R-RRRRRRRRRMhFCR
RRRRRR-R-Rl7FN:HM
RRRRRRRRR--RRRRRRRRpMRHRvBmuXp 
RRRRRRRRR--RRRRRRRR)MRHRvBmuXp 
RRRRRRRRR-- FsssFROM08HH#FM:R
RRRRRR-R-RRRRRRRRRMhFCR
RRRRRR-R-RM)No
C:RRRRRRRR-R-RRRRRR"RR+Z"52#RHR0lNENCl0NHODRD$kFMLkCM88R
RRRRRR-R-R0hFC
#:RRRRRRRR-R-RRRRRRhRRF
MC
RRRRMVkOF0HM+R""RR5pH:RM R)qRp;RRRR)H:RMmRBv upXRR2skC0sBMRmpvu 
X;RRRRRRRR-u-RkFsb#
C:RRRRRRRR-R-RRRRRR)RRCs0kMN#RsEH0lHC0O8RN8HH0FFMRVRRpNRM8)R
RRRRRR-R-RC1bODHNRDPNk:C#
RRRRRRRRR--RRRRRRRRhCFM
RRRRRRRRR--7NFlH
M:RRRRRRRR-R-RRRRRRpRRRRHM)p q
RRRRRRRRR--RRRRRRRR)MRHRvBmuXp 
RRRRRRRRR-- FsssFROM08HH#FM:R
RRRRRR-R-RRRRRRRRRMhFCR
RRRRRR-R-RM)No
C:RRRRRRRR-R-RRRRRR"RR+Z"52#RHR0lNENCl0NHODRD$kFMLkCM88R
RRRRRR-R-R0hFC
#:RRRRRRRR-R-RRRRRRhRRF
MC
RRRRMVkOF0HM+R""RR5pH:RMmRBv upXm_up;q)RR):HBMRmpvu uX_m)pq2R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRCRs0MksRvBmuXp _pumq
);RRRRRRRR-u-RkFsb#
C:RRRRRRRR-R-RRRRRR)RRCs0kMN#RsEH0lHC0O8RN8HH0FFMRVRRpNRM8)R
RRRRRR-R-RC1bODHNRDPNk:C#
RRRRRRRRR--RRRRRRRRhCFM
RRRRRRRRR--7NFlH
M:RRRRRRRR-R-RRRRRRpRRRRHMBumvp_ Xuqmp)MRN83RpqR)t/-=Rv]qa_
uQRRRRRRRR-R-RRRRRR)RRRRHMBumvp_ Xuqmp)MRN83R)qR)t/-=Rv]qa_
uQRRRRRRRR- -RsssFRMOF8HH0F:M#
RRRRRRRRR--RRRRRRRR FsssVRHRqp3)=tRRq-vau]_QR
RRRRRR-R-RRRRRRRRRs sFHsRV3R)qR)t=vR-q_a]uRQ
RRRRR-RR-NR)M:oC
RRRRRRRRR--RRRRRRRRskC#Dv03q>tR=3RjjR
RRRRRR-R-RRRRRRRRRq-vau]_QRR<skC#Dq03)<tR=qRvau]_QR
RRRRRR-R-R0hFC
#:RRRRRRRR-R-RRRRRRhRRF
MC
R
RRkRVMHO0F"MR+5"RRRp:HBMRmpvu RX;RR):H)MR Rqp2RRRR0sCkRsMBumvp; X
RRRRRRRRR--ubksF:#C
RRRRRRRRR--RRRRRRRR)kC0sRM#N0sHE0lCHNOR808HHRFMFpVRR8NMRR)
RRRRR-RR-bR1CNOHDNRPD#kC:R
RRRRRR-R-RRRRRRRRRMhFCR
RRRRRR-R-Rl7FN:HM
RRRRRRRRR--RRRRRRRRpMRHRvBmuXp 
RRRRRRRRR--RRRRRRRR)MRHRq) pR
RRRRRR-R-Rs sFOsRFHM80MHF#R:
RRRRR-RR-RRRRRRRRFRhMRC
RRRRR-RR-NR)M:oC
RRRRRRRRR--RRRRRRRR"5+"ZH2R#NRl0lECNO0HN$DDRLkMF8kMCR8
RRRRR-RR-FRh0:C#
RRRRRRRRR--RRRRRRRRhCFM
R
RRkRVMHO0F"MR+5"RRRp:HBMRmpvu uX_m)pq;)RR:MRHRq) ps2RCs0kMmRBv upXm_up;q)
RRRRRRRRR--ubksF:#C
RRRRRRRRR--RRRRRRRR)kC0sRM#N0sHE0lCHNOR808HHRFMFpVRR8NMRR)
RRRRR-RR-bR1CNOHDNRPD#kC:R
RRRRRR-R-RRRRRRRRRMhFCR
RRRRRR-R-Rl7FN:HM
RRRRRRRRR--RRRRRRRRpMRHRvBmuXp _pumqN)RMp8R3tq)RR/=-avq]Q_u
RRRRRRRRR--RRRRRRRR)MRHRq) pR
RRRRRR-R-Rs sFOsRFHM80MHF#R:
RRRRR-RR-RRRRRRRRsR sRFsHpVR3tq)R-=Rv]qa_
uQRRRRRRRR-)-RNCMo:R
RRRRRR-R-RRRRRRRRR#sCk3D0vRqt>j=R3Rj
RRRRR-RR-RRRRRRRRvR-q_a]u<QRR#sCk3D0qR)t<v=Rq_a]uRQ
RRRRR-RR-FRh0:C#
RRRRRRRRR--RRRRRRRRhCFM
R
RRkRVMHO0F"MR+5"RRRp:H)MR ;qpR:R)RRHMBumvp_ Xuqmp)s2RCs0kMmRBv upXm_up;q)
RRRRRRRRR--ubksF:#C
RRRRRRRRR--RRRRRRRR)kC0sRM#N0sHE0lCHNOR808HHRFMFpVRR8NMRR)
RRRRR-RR-bR1CNOHDNRPD#kC:R
RRRRRR-R-RRRRRRRRRMhFCR
RRRRRR-R-Rl7FN:HM
RRRRRRRRR--RRRRRRRRpMRHRq) pR
RRRRRR-R-RRRRRRRRRH)RMmRBv upXm_upRq)NRM8))3qt=R/Rq-vau]_QR
RRRRRR-R-Rs sFOsRFHM80MHF#R:
RRRRR-RR-RRRRRRRRsR sRFsH)VR3tq)R-=Rv]qa_
uQRRRRRRRR-)-RNCMo:R
RRRRRR-R-RRRRRRRRR#sCk3D0vRqt>j=R3Rj
RRRRR-RR-RRRRRRRRvR-q_a]u<QRR#sCk3D0qR)t<v=Rq_a]uRQ
RRRRR-RR-FRh0:C#
RRRRRRRRR--RRRRRRRRhCFM
R
RRkRVMHO0F"MR-5"RRRp:H)MR ;qpRRRRRR):HBMRmpvu 2XRR0sCkRsMBumvp; X
RRRRRRRRR--ubksF:#C
RRRRRRRRR--RRRRRRRR)kC0sRM#N0sHE0lCH#ORksL0NHO0FFMRVRRplkHM#
R)RRRRRRRR-1-RbHCONPDRNCDk#R:
RRRRR-RR-RRRRRRRRFRhMRC
RRRRR-RR-FR7lMNH:R
RRRRRR-R-RRRRRRRRRHpRM R)qRp
RRRRR-RR-RRRRRRRRRR)HBMRmpvu RX
RRRRR-RR-sR sRFsO8FMHF0HM
#:RRRRRRRR-R-RRRRRRhRRF
MCRRRRRRRR-)-RNCMo:R
RRRRRR-R-RRRRRRRRR""-5RZ2Hl#RNC0ElHN0ODND$MRkLMFk8
C8RRRRRRRR-h-RF#0C:R
RRRRRR-R-RRRRRRRRRMhFCR

RVRRk0MOHRFM"R-"5:RpRRHMBumvp; XR:R)RRHMBumvpR X2CRs0MksRvBmuXp ;R
RRRRRR-R-RsukbCF#:R
RRRRRR-R-RRRRRRRRR0)Ck#sMRHNs0CEl0RHO#0kLs0NOHRFMFpVRRMlHk)#R
RRRRRRRRR--1ObCHRNDPkNDC
#:RRRRRRRR-R-RRRRRRhRRF
MCRRRRRRRR-7-RFHlNMR:
RRRRR-RR-RRRRRRRRRRpHBMRmpvu RX
RRRRR-RR-RRRRRRRRRR)HBMRmpvu RX
RRRRR-RR-sR sRFsO8FMHF0HM
#:RRRRRRRR-R-RRRRRRhRRF
MCRRRRRRRR-)-RNCMo:R
RRRRRR-R-RRRRRRRRR""-5RZ2Hl#RNC0ElHN0ODND$MRkLMFk8
C8RRRRRRRR-h-RF#0C:R
RRRRRR-R-RRRRRRRRRMhFCR

RVRRk0MOHRFM"R-"5:RpRRHMBumvp; XR:R)RRHM)p qRR2RRCRs0MksRvBmuXp ;R
RRRRRR-R-RsukbCF#:R
RRRRRR-R-RRRRRRRRR0)Ck#sMRHNs0CEl0RHO#0kLs0NOHRFMFpVRRMlHk)#R
RRRRRRRRR--1ObCHRNDPkNDC
#:RRRRRRRR-R-RRRRRRhRRF
MCRRRRRRRR-7-RFHlNMR:
RRRRR-RR-RRRRRRRRRRpHBMRmpvu RX
RRRRR-RR-RRRRRRRRRR)H)MR 
qpRRRRRRRR- -RsssFRMOF8HH0F:M#
RRRRRRRRR--RRRRRRRRhCFM
RRRRRRRRR--)oNMCR:
RRRRR-RR-RRRRRRRR-R""25ZRRH#lEN0C0lNHDONDk$RMkLFM88C
RRRRRRRRR--hCF0#R:
RRRRR-RR-RRRRRRRRFRhM
C
RRRRVOkM0MHFR""-Rp5R:MRHRq) pR;R)H:RMmRBv upXm_up2q)R0sCkRsMBumvp_ Xuqmp)R;
RRRRR-RR-kRus#bFCR:
RRRRR-RR-RRRRRRRRCR)0Mks#sRNHl0ECO0HRL#k0OsN0MHFRRFVpHRlMRk#)R
RRRRRR-R-RC1bODHNRDPNk:C#
RRRRRRRRR--RRRRRRRRhCFM
RRRRRRRRR--7NFlH
M:RRRRRRRR-R-RRRRRRpRRRRHM)p q
RRRRRRRRR--RRRRRRRR)MRHRvBmuXp _pumqN)RM)8R3tq)RR/=-avq]Q_u
RRRRRRRRR-- FsssFROM08HH#FM:R
RRRRRR-R-RRRRRRRRRs sFHsRV3R)qR)t=vR-q_a]uRQ
RRRRR-RR-NR)M:oC
RRRRRRRRR--RRRRRRRRskC#Dv03q>tR=3RjjR
RRRRRR-R-RRRRRRRRRq-vau]_QRR<skC#Dq03)<tR=qRvau]_QR
RRRRRR-R-R0hFC
#:RRRRRRRR-R-RRRRRRhRRF
MC
R
RRkRVMHO0F"MR-5"RRRp:HBMRmpvu uX_m)pq;:R)RRHMBumvp_ Xuqmp)R2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRsRRCs0kMmRBv upXm_up;q)
RRRRRRRRR--ubksF:#C
RRRRRRRRR--RRRRRRRR)kC0sRM#N0sHE0lCH#ORksL0NHO0FFMRVRRplkHM#
R)RRRRRRRR-1-RbHCONPDRNCDk#R:
RRRRR-RR-RRRRRRRRFRhMRC
RRRRR-RR-FR7lMNH:R
RRRRRR-R-RRRRRRRRRHpRMmRBv upXm_upRq)NRM8p)3qt=R/Rq-vau]_QR
RRRRRR-R-RRRRRRRRRH)RMmRBv upXm_upRq)NRM8))3qt=R/Rq-vau]_QR
RRRRRR-R-Rs sFOsRFHM80MHF#R:
RRRRR-RR-RRRRRRRRsR sRFsHpVR3tq)R-=Rv]qa_
uQRRRRRRRR-R-RRRRRR RRsssFRRHV))3qtRR=-avq]Q_u
RRRRRRRRR--)oNMCR:
RRRRR-RR-RRRRRRRRCRs#0kD3tvqRR>=j
3jRRRRRRRR-R-RRRRRR-RRv]qa_RuQ<CRs#0kD3tq)RR<=v]qa_
uQRRRRRRRR-h-RF#0C:R
RRRRRR-R-RRRRRRRRRMhFCR

RVRRk0MOHRFM"R-"5:RpRRHMBumvp_ Xuqmp)R;R)H:RM R)qRp2skC0sBMRmpvu uX_m)pq;R
RRRRRR-R-RsukbCF#:R
RRRRRR-R-RRRRRRRRR0)Ck#sMRHNs0CEl0RHO#0kLs0NOHRFMFpVRRMlHk)#R
RRRRRRRRR--1ObCHRNDPkNDC
#:RRRRRRRR-R-RRRRRRhRRF
MCRRRRRRRR-7-RFHlNMR:
RRRRR-RR-RRRRRRRRRRpHBMRmpvu uX_m)pqR8NMRqp3)/tR=vR-q_a]uRQ
RRRRR-RR-RRRRRRRRRR)H)MR 
qpRRRRRRRR- -RsssFRMOF8HH0F:M#
RRRRRRRRR--RRRRRRRR FsssVRHRqp3)=tRRq-vau]_QR
RRRRRR-R-RM)No
C:RRRRRRRR-R-RRRRRRsRRCD#k0q3vt=R>Rjj3
RRRRRRRRR--RRRRRRRR-avq]Q_uRs<RCD#k0)3qt=R<Ravq]Q_u
RRRRRRRRR--hCF0#R:
RRRRR-RR-RRRRRRRRFRhM
C
RRRRVOkM0MHFR""*Rp5R:MRHRvBmuXp ;)RR:MRHRvBmuXp Rs2RCs0kMmRBv upXR;
RRRRR-RR-kRus#bFCR:
RRRRR-RR-RRRRRRRRCR)0Mks#sRNHl0ECO0HRDlk0DHbH0ONHRFMFpVRR8NMRR)
RRRRR-RR-bR1CNOHDNRPD#kC:R
RRRRRR-R-RRRRRRRRRMhFCR
RRRRRR-R-Rl7FN:HM
RRRRRRRRR--RRRRRRRRpMRHRvBmuXp 
RRRRRRRRR--RRRRRRRR)MRHRvBmuXp 
RRRRRRRRR-- FsssFROM08HH#FM:R
RRRRRR-R-RRRRRRRRRMhFCR
RRRRRR-R-RM)No
C:RRRRRRRR-R-RRRRRR"RR*Z"52#RHR0lNENCl0NHODRD$kFMLkCM88R
RRRRRR-R-R0hFC
#:RRRRRRRR-R-RRRRRRhRRF
MC
RRRRMVkOF0HM*R""RR5pH:RMmRBv upXR;R)H:RM R)q2pRRCRs0MksRvBmuXp ;R
RRRRRR-R-RsukbCF#:R
RRRRRR-R-RRRRRRRRR0)Ck#sMRHNs0CEl0RHOl0kDHHbDOHN0FFMRVRRpNRM8)R
RRRRRR-R-RC1bODHNRDPNk:C#
RRRRRRRRR--RRRRRRRRhCFM
RRRRRRRRR--7NFlH
M:RRRRRRRR-R-RRRRRRpRRRRHMBumvp
 XRRRRRRRR-R-RRRRRR)RRRRHM)p q
RRRRRRRRR-- FsssFROM08HH#FM:R
RRRRRR-R-RRRRRRRRRMhFCR

RRRRR-RR-NR)M:oC
RRRRRRRRR--RRRRRRRR"5*"ZH2R#NRl0lECNO0HN$DDRLkMF8kMCR8
RRRRR-RR-FRh0:C#
RRRRRRRRR--RRRRRRRRhCFM
R
RRkRVMHO0F"MR*5"RRRp:H)MR ;qpR:R)RRHMBumvpR X2CRs0MksRvBmuXp ;R
RRRRRR-R-RsukbCF#:R
RRRRRR-R-RRRRRRRRR0)Ck#sMRHNs0CEl0RHOl0kDHHbDOHN0FFMRVRRpNRM8)R
RRRRRR-R-RC1bODHNRDPNk:C#
RRRRRRRRR--RRRRRRRRhCFM
RRRRRRRRR--7NFlH
M:RRRRRRRR-R-RRRRRRpRRRRHM)p q
RRRRRRRRR--RRRRRRRR)MRHRvBmuXp 
RRRRRRRRR-- FsssFROM08HH#FM:R
RRRRRR-R-RRRRRRRRRMhFCR
RRRRRR-R-RM)No
C:RRRRRRRR-R-RRRRRR"RR*Z"52#RHR0lNENCl0NHODRD$kFMLkCM88R
RRRRRR-R-R0hFC
#:RRRRRRRR-R-RRRRRRhRRF
MC
RRRRMVkOF0HM*R""RR5pH:RMmRBv upXm_up;q)RR):HBMRmpvu uX_m)pq2R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRCRs0MksRvBmuXp _pumq
);RRRRRRRR-u-RkFsb#
C:RRRRRRRR-R-RRRRRR)RRCs0kMN#RsEH0lHC0OkRlDb0HDNHO0MHFRRFVpMRN8
R)RRRRRRRR-1-RbHCONPDRNCDk#R:
RRRRR-RR-RRRRRRRRFRhMRC
RRRRR-RR-FR7lMNH:R
RRRRRR-R-RRRRRRRRRHpRMmRBv upXm_upRq)NRM8p)3qt=R/Rq-vau]_QR
RRRRRR-R-RRRRRRRRRH)RMmRBv upXm_upRq)NRM8))3qt=R/Rq-vau]_QR
RRRRRR-R-Rs sFOsRFHM80MHF#R:
RRRRR-RR-RRRRRRRRsR sRFsHpVR3tq)R-=Rv]qa_
uQRRRRRRRR-R-RRRRRR RRsssFRRHV))3qtRR=-avq]Q_u
RRRRRRRRR--)oNMCR:
RRRRR-RR-RRRRRRRRCRs#0kD3tvqRR>=j
3jRRRRRRRR-R-RRRRRR-RRv]qa_RuQ<CRs#0kD3tq)RR<=v]qa_
uQRRRRRRRR-h-RF#0C:R
RRRRRR-R-RRRRRRRRRMhFCR

RVRRk0MOHRFM"R*"5:RpRRHM)p q;)RR:MRHRvBmuXp _pumqR)2skC0sBMRmpvu uX_m)pq;R
RRRRRR-R-RsukbCF#:R
RRRRRR-R-RRRRRRRRR0)Ck#sMRHNs0CEl0RHOl0kDHHbDOHN0FFMRVRRpNRM8)R
RRRRRR-R-RC1bODHNRDPNk:C#
RRRRRRRRR--RRRRRRRRhCFM
RRRRRRRRR--7NFlH
M:RRRRRRRR-R-RRRRRRpRRRRHM)p q
RRRRRRRRR--RRRRRRRR)MRHRvBmuXp _pumqN)RM)8R3tq)RR/=-avq]Q_u
RRRRRRRRR-- FsssFROM08HH#FM:R
RRRRRR-R-RRRRRRRRRs sFHsRV3R)qR)t=vR-q_a]uRQ
RRRRR-RR-NR)M:oC
RRRRRRRRR--RRRRRRRRskC#Dv03q>tR=3RjjR
RRRRRR-R-RRRRRRRRRq-vau]_QRR<skC#Dq03)<tR=qRvau]_QR
RRRRRR-R-R0hFC
#:RRRRRRRR-R-RRRRRRhRRF
MC
RRRRMVkOF0HM*R""RR5pH:RMmRBv upXm_up;q)R:R)RRHM)p q2CRs0MksRvBmuXp _pumq
);RRRRRRRR-u-RkFsb#
C:RRRRRRRR-R-RRRRRR)RRCs0kMN#RsEH0lHC0OkRlDb0HDNHO0MHFRRFVpMRN8
R)RRRRRRRR-1-RbHCONPDRNCDk#R:
RRRRR-RR-RRRRRRRRFRhMRC
RRRRR-RR-FR7lMNH:R
RRRRRR-R-RRRRRRRRRHpRMmRBv upXm_upRq)NRM8p)3qt=R/Rq-vau]_QR
RRRRRR-R-RRRRRRRRRH)RM R)qRp
RRRRR-RR-sR sRFsO8FMHF0HM
#:RRRRRRRR-R-RRRRRR RRsssFRRHVp)3qtRR=-avq]Q_u
RRRRRRRRR--)oNMCR:
RRRRR-RR-RRRRRRRRCRs#0kD3tvqRR>=j
3jRRRRRRRR-R-RRRRRR-RRv]qa_RuQ<CRs#0kD3tq)RR<=v]qa_
uQRRRRRRRR-h-RF#0C:R
RRRRRR-R-RRRRRRRRRMhFC


RRRRVOkM0MHFR""/Rp5R:MRHRq) pR;R)H:RMmRBv upXRR2skC0sBMRmpvu 
X;RRRRRRRR-u-RkFsb#
C:RRRRRRRR-R-RRRRRR)RRCs0kMN#RsEH0lHC0OHR8PHH#FFMRVRRpL)$R
RRRRRRRRR--1ObCHRNDPkNDC
#:RRRRRRRR-R-RRRRRRhRRF
MCRRRRRRRR-7-RFHlNMR:
RRRRR-RR-RRRRRRRRRRpH)MR 
qpRRRRRRRR-R-RRRRRR)RRRRHMBumvpR XNRM8)=R/Ravq]Z_B 
)mRRRRRRRR- -RsssFRMOF8HH0F:M#
RRRRRRRRR--RRRRRRRR FsssVRHR=)RRavq]Z_B 
)mRRRRRRRR-)-RNCMo:R
RRRRRR-R-RRRRRRRRR""/5RZ2Hl#RNC0ElHN0ODND$MRkLMFk8
C8RRRRRRRR-h-RF#0C:R
RRRRRR-R-RRRRRRRRRMhFCR

RVRRk0MOHRFM"R/"5:RpRRHMBumvp; XR:R)RRHMBumvpR X2CRs0MksRvBmuXp ;R
RRRRRR-R-RsukbCF#:R
RRRRRR-R-RRRRRRRRR0)Ck#sMRHNs0CEl0RHO8HHP#MHFRRFVp$RLRR)
RRRRR-RR-bR1CNOHDNRPD#kC:R
RRRRRR-R-RRRRRRRRRMhFCR
RRRRRR-R-Rl7FN:HM
RRRRRRRRR--RRRRRRRRpMRHRvBmuXp 
RRRRRRRRR--RRRRRRRR)MRHRvBmuXp R8NMR/)R=qRvaB]_Zm )
RRRRRRRRR-- FsssFROM08HH#FM:R
RRRRRR-R-RRRRRRRRRs sFHsRVRR)=qRvaB]_Zm )
RRRRRRRRR--)oNMCR:
RRRRR-RR-RRRRRRRR/R""25ZRRH#lEN0C0lNHDONDk$RMkLFM88C
RRRRRRRRR--hCF0#R:
RRRRR-RR-RRRRRRRRFRhM
C
RRRRVOkM0MHFR""/Rp5R:MRHRvBmuXp ;)RR:MRHRq) pRR2RsRRCs0kMmRBv upXR;
RRRRR-RR-kRus#bFCR:
RRRRR-RR-RRRRRRRRCR)0Mks#sRNHl0ECO0HRP8HHF#HMVRFRLpR$
R)RRRRRRRR-1-RbHCONPDRNCDk#R:
RRRRR-RR-RRRRRRRRFRhMRC
RRRRR-RR-FR7lMNH:R
RRRRRR-R-RRRRRRRRRHpRMmRBv upXR
RRRRRR-R-RRRRRRRRRH)RM R)qNpRM)8RRR/=j
3jRRRRRRRR- -RsssFRMOF8HH0F:M#
RRRRRRRRR--RRRRRRRR FsssVRHR=)RRjj3
RRRRRRRRR--)oNMCR:
RRRRR-RR-RRRRRRRR/R""25ZRRH#lEN0C0lNHDONDk$RMkLFM88C
RRRRRRRRR--hCF0#R:
RRRRR-RR-RRRRRRRRFRhM
C
RRRRVOkM0MHFR""/Rp5R:MRHRvBmuXp _pumqR);)H:RMmRBv upXm_up2q)
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR0sCkRsMBumvp_ Xuqmp)R;
RRRRR-RR-kRus#bFCR:
RRRRR-RR-RRRRRRRRCR)0Mks#sRNHl0ECO0HRP8HHF#HMVRFRLpR$
R)RRRRRRRR-1-RbHCONPDRNCDk#R:
RRRRR-RR-RRRRRRRRFRhMRC
RRRRR-RR-FR7lMNH:R
RRRRRR-R-RRRRRRRRRHpRMmRBv upXm_upRq)NRM8p)3qt=R/Rq-vau]_QR
RRRRRR-R-RRRRRRRRRH)RMmRBv upXm_upRq)NRM8))3qt=R/Rq-vau]_QR
RRRRRR-R-RRRRRRRRRv)3q>tRRjj3
RRRRRRRRR-- FsssFROM08HH#FM:R
RRRRRR-R-RRRRRRRRRs sFHsRV3R)vRqt<j=R3Rj
RRRRR-RR-RRRRRRRRsR sRFsHpVR3tq)R-=Rv]qa_
uQRRRRRRRR-R-RRRRRR RRsssFRRHV))3qtRR=-avq]Q_u
RRRRRRRRR--)oNMCR:
RRRRR-RR-RRRRRRRRCRs#0kD3tvqRR>=j
3jRRRRRRRR-R-RRRRRR-RRv]qa_RuQ<CRs#0kD3tq)RR<=v]qa_
uQRRRRRRRR-h-RF#0C:R
RRRRRR-R-RRRRRRRRRMhFCR

RVRRk0MOHRFM"R/"5:RpRRHM)p q;)RR:MRHRvBmuXp _pumqR)2skC0sBMRmpvu uX_m)pq;R
RRRRRR-R-RsukbCF#:R
RRRRRR-R-RRRRRRRRR0)Ck#sMRHNs0CEl0RHO8HHP#MHFRRFVp$RLRR)
RRRRR-RR-bR1CNOHDNRPD#kC:R
RRRRRR-R-RRRRRRRRRMhFCR
RRRRRR-R-Rl7FN:HM
RRRRRRRRR--RRRRRRRRpMRHRq) pR
RRRRRR-R-RRRRRRRRRH)RMmRBv upXm_upRq)NRM8))3qt=R/Rq-vau]_QR
RRRRRR-R-RRRRRRRRRv)3q>tRRjj3
RRRRRRRRR-- FsssFROM08HH#FM:R
RRRRRR-R-RRRRRRRRRs sFHsRV3R)vRqt<j=R3Rj
RRRRR-RR-RRRRRRRRsR sRFsH)VR3tq)R-=Rv]qa_
uQRRRRRRRR-)-RNCMo:R
RRRRRR-R-RRRRRRRRR#sCk3D0vRqt>j=R3Rj
RRRRR-RR-RRRRRRRRvR-q_a]u<QRR#sCk3D0qR)t<v=Rq_a]uRQ
RRRRR-RR-FRh0:C#
RRRRRRRRR--RRRRRRRRhCFM
R
RRkRVMHO0F"MR/5"RRRp:HBMRmpvu uX_m)pq;)RR:MRHRq) ps2RCs0kMmRBv upXm_up;q)
RRRRRRRRR--ubksF:#C
RRRRRRRRR--RRRRRRRR)kC0sRM#N0sHE0lCH8ORH#PHHRFMFpVRRRL$)R
RRRRRR-R-RC1bODHNRDPNk:C#
RRRRRRRRR--RRRRRRRRhCFM
RRRRRRRRR--7NFlH
M:RRRRRRRR-R-RRRRRRpRRRRHMBumvp_ Xuqmp)MRN83RpqR)t/-=Rv]qa_
uQRRRRRRRR-R-RRRRRR)RRRR/=j
3jRRRRRRRR- -RsssFRMOF8HH0F:M#
RRRRRRRRR--RRRRRRRR FsssVRHRqp3)=tRRq-vau]_QR
RRRRRR-R-RRRRRRRRRs sFHsRVRR)=3RjjR
RRRRRR-R-RM)No
C:RRRRRRRR-R-RRRRRRsRRCD#k0q3vt=R>Rjj3
RRRRRRRRR--RRRRRRRR-avq]Q_uRs<RCD#k0)3qt=R<Ravq]Q_u
RRRRRRRRR--hCF0#R:
RRRRR-RR-RRRRRRRRFRhMCC
MR8Rv]qa_vBmuXp ;-
------------------------------------------------------------------------
--
-RbBF$osHE40RgRgnLQ$R 3  RDqDRosHER0#sCC#s8PC3-
-
R--a#EHRk#FsROCVCHDRRH#NHMRMsVFlHN0PbCRNRs0FQVR R  1R084nj(34.-g,gnR Q  0R1NNM8s
8R-e-R]R7pvEN0C0lNHDONROuN	CNo#a3RERH##sFkOVCRHRDClRN$MRF0LOCRFCbH8#,RF,D8RRFs
R--HDMOk88CR0IHEFR#VN0Is0CRERN0H##RFRD8IEH0FRk0I0sH0RCMblCsHH##FVMRsRFl0RECQ   
R--1M0N88Ns#CR7b0Nsl0CM3ERaH##RFOksCHRVDlCRNL$RC#RkC08RFlRHblDCCRM00#EHRN#0Ms8N8-R
-MRN8NRl$CRLR#8H0LsHk80CRRHMObFlH8DCRsVFlMRHR$NMRMlNMRCs#DFRFRMoN0#RE
CR-O-RFHlbDRC8VlFsRC8F#FRM0DRNDRFI8CHsO80RClOFbNHD0MHFRRFV0RECFosHHDMNRk#FsROCVCHD3-
-RHaE#FR#kCsORDVHCNRl$CRLRbOFHRC8VRFsHHM8PkH8NkDR#LCRCC0ICDMRHMOC#RC8ks#C#
3R-a-RERH##sFkOVCRHRDCHb#RsHFP8RC8FNMRM1RqRRQ1LHN##a3REQCR R  8OH#DlNH#hRqY-R
-qRW)h)qa YRX u)1m1R)vRQu pQ7hRQB7pzQRhtqRhYW)q)qYhaRRmwvB )]aqhqpAQQRaY
R--qRh7whQa R11wRm)zR1 wRm)qqRu)BaQz)pqR)uzu m13ERaC#RkCFsRVER0CFR#kCsOR-
-RDVHCER#NRDDHCM8lVMH$MRN8FREDQ8R R  ElNsD#C#RFVslMRN$NR8lCNo#sRFRNDHLHHD0
$R-N-RsHH#MFoRkF0RVER0C#RkCER0CFsCV-3
--
-R0aHDRC:RRRRR0R1NNM8se8R]R7pvEN0C0lNHDONROuN	CNo#QR5 R  1R084nj(34.-g,gn
R--RRRRRRRRRRRRRavq]m_Bv upX-2
--
-RLpHs$Ns:RRRRERaHb#RNNO	o#CREDNDRRLCObFlH8DCR0HMFRRNDsHLN
s$-R-RRRRRRRRRRRRR#L$lFODHN$DDRlMNCQ8R 3  

---7-RCDPCFsbC#R:RQ   R17qB]Re7vpRNC0ElHN0ORNDu	NON#oCRsWF	oHMRFtsk-b
--
-RsukbCF#:RRRRERaHb#RNNO	oLCRFR8$HN#RRMMFMlFsNP0HClRHblDCCNM00MHFRRFV0REC
R--RRRRRRRRRRRRRMVkOF0HMHND08$RCMVHCH8RMER0CqRvaB]_mpvu bXRNNO	o8CRCNODsHN0F
M3---
-HRplNH00MHF:aRREPCRNCDk#CRoMNCs0RC8L0$REVCRk0MOH#FMRRHM0#EHRObN	CNoR$lN
R--RRRRRRRRRRRRRsPN$sRVFblRDVN0FRsl0bFRDVN0F,slR8NMRC0ERCbsOHH#FFMRVCRs#0kD#-
-RRRRRRRRRRRRR#RHRDFM$kRoNMsN08CCRR0FL0CRElCRHlMHkslRCHJksRC8LQ$R R  1R084nj(
R--RRRRRRRRRRRRRg-4g
d3---
-FRh0:C#
R--RRRRRRRRRRRRRCaERN"bOo	NCCR8OsDNNF0HM8"RCMVHC0#RE0CR$#bC,kR#Lb0$CR#,N
M8-R-RRRRRRRRRRRRR8DCON0sNH#FMRRFVv]qa_vBmuXp 3-
-RRRRRRRRRRRRRERaC0R#NNM8sl8RNC0ElHN0ORND8HCVMHH0FNMRMO8RFCMPMF0HMRNDlMCNH
Mo-R-RRRRRRRRRRRRRF0VRElCRNC0ElHN0ORNDVOkM0MHF#ER0NN0RsbCRNRs0F0VRERH##M0N88Ns
R--RRRRRRRRRRRRRbsCsCC#M00REVCRFNslDCR#l0NMHRO#F0VREHCRlCbDl0CMNF0HMVRFRC0E
R--RRRRRRRRRRRRRavq]m_Bv upXNRbOo	NCCR8OsDNNF0HMR3RaRECbbksFR#CF0VRE-C
-RRRRRRRRRRRRvRRq_a]BumvpR Xb	NONRoCL$F8RRH#0OFRDHNsV#$RkROE#NClMO0H#MRN8-
-RRRRRRRRRRRRRsRbF8PHCRRNo8kHCMDHCFRVslRHblDCCNM00MHF#FR0RsPCHRV$0HECs-
-RRRRRRRRRRRRRlRHblDCCNM00MHFRRFVv]qa_vBmuXp 3aRRFRFD8CCPDCFbsl#RNO$RE#FFCFR0
R--RRRRRRRRRRRRRbHlDCClM00REbCRNNO	oLCRFR8$H0MRElCRFR#0CHVVOMHC0NRlMsMC
R--RRRRRRRRRRRRRNNPHLDND0CRFER0C
l3---
--R--------------------------------------------------------------------------
---e-RCHs#FRMRRRR:4
36-7-RNR0CRRRRRRR:.KcRkRD$4ngg
R-------------------------------------------------------------------------------k

#WCRm3)iv]qa_q) pD3ND
;
b	NONRoCL$F8Ravq]m_Bv upX#RH
R
RR-R-
RRRRR-- NJkD$H0R8NMRCQMJDkNHR0$msbCNs0F#FRVsmRBv upXm_up
q)RRRR-R-
RVRRk0MOHRFM"R="5:RpRRHMBumvp_ Xuqmp)R;R)H:RMmRBv upXm_upRq)2CRs0MksRmAmph q
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR#RH
RRRRRRRRR--7OC#s0HbH:FM
RRRRRRRRR--RRRRR1RRCVCRk0MOHRFM8DCON0sNHRFMHQMR R  1R084nj(34.-g
gnRRRRRRRR-h-RF#0C:R
RRRRRR-R-RRRRRRRRN)2RCs0kMw#Rq p1RRFMCFsssR
RRCRLo
HMRRRRRRRR-B-RE	CORDPNH08H$VRFRbHMkN0RslokC#M0
RRRRRRRRRHV53RpqR)t=vR-q_a]u2QRRC0EMR
RRRRRRRRRRRRRR#RN#0CsRpwq1R 
RRRRRRRRRRRRRRRRRRRRRRRRRsRRCsbF0pR"3tq)R-=Rv]qa_RuQH=MR5)p,2R"
RRRRRRRRRRRRRRRRRRRRRRRRR#RRCsPCHR0$ m)))R;
RRRRRRRRRRRRRsRRCs0kMqRwp;1 
RRRRRRRR8CMR;HV
R
RRRRRRVRHR)5R3tq)R-=Rv]qa_RuQ2ER0CRM
RRRRRRRRRRRRRNRR#s#C0qRwp
1 RRRRRRRRRRRRRRRRRRRRRRRRRRRRsFCbs"0R))3qtRR=-avq]Q_uRRHM=,5p)
2"RRRRRRRRRRRRRRRRRRRRRRRRRRRR#CCPs$H0R) )m
);RRRRRRRRRRRRRRRRskC0swMRq p1;R
RRRRRRMRC8VRH;R

RRRRR-RR-CRt0bR#CNOHDNRPD#kC
RRRRRRRRRHV53RpvRqt=3RjjMRN83R)vRqt=3RjjRR20MEC
RRRRRRRRRRRRRRRR0sCkRsMa )z;R
RRRRRRMRC8VRH;R

RRRRR-RR-CRt0NRPDRkCVRFsoCCMsRNDOCN#
RRRRRRRRRHV53RpvRqt=3R)vRqtNRM8p)3qtRR=))3qtRR20MEC
RRRRRRRRRRRRRRRR0sCkRsMa )z;R
RRRRRRMRC8VRH;R

RRRRRsRRCs0kMqRwp;1 
RRRR8CMR""=;


RRRRVOkM0MHFR="/"RR5pH:RMmRBv upXm_up;q)R:R)RRHMBumvp_ Xuqmp)RR2skC0sAMRm mpqRh
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRHR#
RRRRR-RR-CR7#HOsbF0HMR:
RRRRR-RR-RRRRRRRRC1CRMVkOF0HMCR8OsDNNF0HMMRHR Q  0R18jR4(.n3-g4gnR
RRRRRR-R-R0hFC
#:RRRRRRRR-R-RRRRRR2RNR0)Ck#sMRpwq1F RMsRCs
FsRRRRLHCoMR
RRRRRR-R-RCBEOP	RN8DHHR0$FHVRM0bkRoNskMlC0R#
RRRRRHRRVRR5p)3qtRR=-avq]Q_uR02RE
CMRRRRRRRRRRRRRRRRNC##sw0Rq p1
RRRRRRRRRRRRRRRRRRRRRRRRRRRRbsCFRs0"qp3)=tRRq-vau]_QMRHR5/=p2,)"R
RRRRRRRRRRRRRRRRRRRRRRRRRRCR#PHCs0 $R)))m;R
RRRRRRRRRRRRRRCRs0MksRpwq1
 ;RRRRRRRRCRM8H
V;
RRRRRRRRRHV53R)qR)t=vR-q_a]u2QRRC0EMR
RRRRRRRRRRRRRR#RN#0CsRpwq1R 
RRRRRRRRRRRRRRRRRRRRRRRRRsRRCsbF0)R"3tq)R-=Rv]qa_RuQH/MR=,5p)
2"RRRRRRRRRRRRRRRRRRRRRRRRRRRR#CCPs$H0R) )m
);RRRRRRRRRRRRRRRRskC0swMRq p1;R
RRRRRRMRC8VRH;R

RRRRR-RR-CRt0bR#CNOHDNRPD#kC
RRRRRRRRRHV53RpvRqt=3RjjMRN83R)vRqt=3RjjRR20MEC
RRRRRRRRRRRRRRRR0sCkRsMw1qp R;
RRRRRCRRMH8RV
;
RRRRRRRR-t-RCP0RNCDkRsVFRMoCCDsNR#ONCR
RRRRRRVRHRp5R3tvqR)=R3tvqR8NMRqp3)=tRRq)3)2tRRC0EMR
RRRRRRRRRRRRRRCRs0MksRpwq1
 ;RRRRRRRRCRM8H
V;
RRRRRRRR0sCkRsMa )z;R
RRMRC8/R"=
";
RRRR
--RRRR-m-R0sECRMwkOF0HM1#R00NsRs]CCR
RR-R-
R
RRkRVMHO0FtMR ua_)BQhQpuq_peqzX 5:MRHRq) pRR2skC0suMR)BQhQpuq_peqzH R#R
RRRRRR-R-R#7CObsH0MHF:R
RRRRRR-R-RRRRRRRR1RCCVOkM0MHFRO8CDNNs0MHFRRHMQ   R810R(4jn-3.4ngg
RRRRRRRRR--hCF0#R:
RRRRR-RR-RRRRRRRRMhFCR
RRRRRRNRPsLHNDaCR :vuRq) pR;
RLRRCMoH
RRRRRRRRR--BOEC	VRHRsNDC$N8RbNRsOHMHDbNRDPNkRC
RRRRRHRRVRR5XRR>-avq]Q_uR8NMR<XR=qRvau]_QRR20MEC
RRRRRRRRRRRRRRRR0sCkRsMuh)QBqQupq_ep'z 5;X2
RRRRRRRR8CMR;HV
R
RRRRRR-R-R0tCRHbsMbOHNPDRNCDk
RRRRRRRRva u=R:R
X;RRRRRRRRIDEHCRR5au vRR<=-avq]Q_uRD2RF
FbRRRRRRRRRRRRRRRRau vRR:=au vRv+Rq_a].Q_u;R
RRRRRRMRC8FRDF
b;RRRRRRRRIDEHCaR5 Rvu>qRvau]_QRR2DbFF
RRRRRRRRRRRRRRRRva u=R:Rva uRR-v]qa_u._QR;
RRRRRCRRMD8RF;Fb
R
RRRRRRCRs0MksRQu)huBQqep_q pz' 5av;u2
RRRR8CMRat _Qu)huBQqep_q pz;R

RVRRk0MOHRFMBpvuX:5XRRHM)p q;YRR:MRHRq) p=R:Rjj3Rs2RCs0kMmRBv upX#RH
RRRRRRRRR--7OC#s0HbH:FM
RRRRRRRRR--RRRRR1RRCVCRk0MOHRFM8DCON0sNHRFMHQMR R  1R084nj(34.-g
gnRRRRRRRR-h-RF#0C:R
RRRRRR-R-RRRRRRRRhCFM
RRRRoLCHRM
RRRRRsRRCs0kMmRBv upXX'5,2RY;R
RRMRC8vRBu;pX
R
RRkRVMHO0FuMRm)pq__amBumvp5 XZH:RMmRBv upXm_upRq)2CRs0MksRvBmuXp R
H#RRRRRRRR-7-RCs#OHHb0F
M:RRRRRRRR-R-RRRRRRCR1CkRVMHO0F8MRCNODsHN0FHMRM RQ 1 R048Rj3(n.g-4gRn
RRRRR-RR-FRh0:C#
RRRRRRRRR--RRRRRNRR2CR)0Mks#qRvaB]_Zm )RRFMCFsssR
RRCRLo
HMRRRRRRRR-B-RE	CORDPNH08H$VRFRbHMkN0RslokC#M0
RRRRRRRRRHV53RZqR)t=vR-q_a]u2QRRC0EMR
RRRRRRRRRRRRRR#RN#0CsRpwq1R 
RRRRRRRRRRRRRRRRRRRRRCRsb0FsR3"ZqR)t=vR-q_a]uHQRMmRup_q)aBm_mpvu ZX52R"
RRRRRRRRRRRRRRRRRRRRRCR#PHCs0 $R)))m;R
RRRRRRRRRRRRRRCRs0MksRavq]Z_B ;)m
RRRRRRRR8CMR;HV
R
RRRRRR-R-R0tCRDPNkVCRFosRCsMCNODRN
#CRRRRRRRRskC0sBMRmpvu 5X'RvZ3qBt*mZ153tq)2Z,R3tvq*h1Q5qZ3)Rt22R;
RCRRMu8Rm)pq__amBumvp; X



RRRRVOkM0MHFRvBmuXp __amuqmp):5ZRRHMBumvpR X2CRs0MksRvBmuXp _pumqH)R#R
RRRRRR-R-R#7CObsH0MHF:R
RRRRRR-R-RRRRRRRR1RCCVOkM0MHFRO8CDNNs0MHFRRHMQ   R810R(4jn-3.4ngg
RRRRRRRRR--hCF0#R:
RRRRR-RR-RRRRRRRRMhFCR
RRRRRRNRPsLHNDaCR :vuRq) pR;
RLRRCMoH
RRRRRRRRR--tRC0PkNDCFRVsbR#CNOHDNRO#
C#RRRRRRRRH5VRR)Z3 RR=jR3j2ER0CRM
RRRRRRRRRHRRVRR5Zv3QRj=R32jRRC0EMR
RRRRRRRRRRRRRRCRs0MksRvBmuXp _pumq5)'j,3jRjj32R;
RRRRRRRRRCRRDV#HRZ5R3RQv>3RjjRR20MEC
RRRRRRRRRRRRRRRR0sCkRsMBumvp_ Xuqmp)Z'53,QvRavq]Q_u_ me)2_.;R
RRRRRRRRRRDRC#RC
RRRRRRRRRRRRRsRRCs0kMmRBv upXm_up'q)53-ZQRv,-avq]Q_u_ me)2_.;R
RRRRRRRRRRMRC8VRH;R
RRRRRRMRC8VRH;R

RRRRRHRRVRR5Zv3QRj=R32jRRC0EMR
RRRRRRRRRRVRHRZ5R3R) =3RjjRR20MEC
RRRRRRRRRRRRRRRR0sCkRsMBumvp_ Xuqmp)j'53Rj,j23j;R
RRRRRRRRRRDRC#RHV53RZ)> RRjj3R02RE
CMRRRRRRRRRRRRRRRRskC0sBMRmpvu uX_m)pq'35Z)R ,j23j;R
RRRRRRRRRRDRC#RC
RRRRRRRRRRRRRsRRCs0kMmRBv upXm_up'q)53-Z)R ,v]qa_2uQ;R
RRRRRRRRRRMRC8VRH;R
RRRRRRMRC8VRH;R

RRRRR-RR-CRt0sRbHHMObRNDPkNDCFRVsCRoMNCsDNRO#RC
RRRRRaRR Rvu:q=R)qBah35ZQRv,Z 3)2
;
RRRRRRRRskC0sBMRmpvu uX_m)pq'T51)Za53*) Z 3)RZ+R3*QvZv3Q2R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRt_ auh)QBqQupq_ep5z au v2
2;RRRRCRM8Bumvp_ Xaum_m)pq;R

RVRRk0MOHRFM"1qA":5ZRRHMBumvpR X2CRs0MksR1umQeaQ  _)qHpR#R
RRRRRR-R-R#7CObsH0MHF:R
RRRRRR-R-RRRRRRRR1RCCVOkM0MHFRO8CDNNs0MHFRRHMQ   R810R(4jn-3.4ngg
RRRRRRRRR--hCF0#R:
RRRRR-RR-RRRRRRRRRN2q5A1Z=2RR)1Ta35Z)Z *3R) +3RZQZv*32Qv
R
RRCRLo
HMRRRRRRRR-t-RCP0RNCDkRsVFRMoCCDsNR#ONCR
RRRRRRCRs0MksR1umQeaQ  _)q5p'1aT)5)Z3 3*Z)+ RRQZ3v3*ZQ2v2;R
RRMRC8qR"A;1"
R
RRkRVMHO0F"MRq"A15RZ:HBMRmpvu uX_m)pqRs2RCs0kMmRu1QQae) _ RqpHR#
RRRRR-RR-CR7#HOsbF0HMR:
RRRRR-RR-RRRRRRRRC1CRMVkOF0HMCR8OsDNNF0HMMRHR Q  0R18jR4(.n3-g4gnR
RRRRRR-R-R0hFC
#:RRRRRRRR-R-RRRRRR2RNR1qA5RZ2=3RZv
qtRRRRRRRR-R-RRRRRR2RLR0)Ck#sMRjj3RRFMCFsssR

RLRRCMoH
RRRRRRRRR--BOEC	NRPDHH80F$RVMRHbRk0Nksol0CM#R
RRRRRRVRHRZ5R3tq)R-=Rv]qa_RuQ2ER0CRM
RRRRRRRRRRRRRRRRR#N#CRs0w1qp R
RRRRRRRRRRRRRRRRRRRRRRRRRRCRsb0FsR3"ZqR)t=vR-q_a]uHQRMARq125Z"R
RRRRRRRRRRRRRRRRRRRRRRRRRRCR#PHCs0 $R)))m;R
RRRRRRRRRRRRRRRRRskC0sjMR3
j;RRRRRRRRCRM8H
V;
RRRRRRRRR--tRC0PkNDCFRVsCRoMNCsDNRO#RC
RRRRRsRRCs0kM3RZv;qt
RRRR8CMRA"q1
";
R
RRkRVMHO0FqMR)Zt5:MRHRvBmuXp Rs2RCs0kM)RuQQhBu_qpezqp #RH
RRRRRRRRR--7OC#s0HbH:FM
RRRRRRRRR--RRRRR1RRCVCRk0MOHRFM8DCON0sNHRFMHQMR R  1R084nj(34.-g
gnRRRRRRRR-h-RF#0C:R
RRRRRR-R-RRRRRRRRNq2R)Zt52RR=qa)BqZh53,QvR)Z3 
2
RRRRRRRRPHNsNCLDR Zav:uRRvBmuXp _pumq
);RRRRLHCoMR
RRRRRR-R-R0tCRDPNkVCRFosRCsMCNODRN
#CRRRRRRRRZva u=R:RvBmuXp __amuqmp)25Z;R
RRRRRRCRs0MksR Zavqu3)
t;RRRRCRM8q;)t
R
RRkRVMHO0FqMR)Zt5:MRHRvBmuXp _pumq2)RR0sCkRsMuh)QBqQupq_epRz HR#
RRRRR-RR-CR7#HOsbF0HMR:
RRRRR-RR-RRRRRRRRC1CRMVkOF0HMCR8OsDNNF0HMMRHR Q  0R18jR4(.n3-g4gnR
RRRRRR-R-R0hFC
#:RRRRRRRR-R-RRRRRR2RNRtq)5RZ2=3RZq
)tRRRRRRRR-R-RRRRRR2RLR0)Ck#sMRjj3RRFMCFsssR

RLRRCMoH
RRRRRRRRR--BOEC	NRPDHH80F$RVMRHbRk0Nksol0CM#R
RRRRRRVRHRZ5R3tq)R-=Rv]qa_RuQ2ER0CRM
RRRRRRRRRRRRRRRRR#N#CRs0w1qp R
RRRRRRRRRRRRRRRRRRRRRRRRRRCRsb0FsR3"ZqR)t=vR-q_a]uHQRM)Rqt25Z"R
RRRRRRRRRRRRRRRRRRRRRRRRRRCR#PHCs0 $R)))m;R
RRRRRRRRRRRRRRRRRskC0sjMR3
j;RRRRRRRRCRM8H
V;
RRRRRRRRR--tRC0PkNDCFRVsCRoMNCsDNRO#RC
RRRRRsRRCs0kM3RZq;)t
RRRR8CMRtq);R

RVRRk0MOHRFM"R-"5RZ:HBMRmpvu 2XRR0sCkRsMBumvpR XHR#
RRRRR-RR-CR7#HOsbF0HMR:
RRRRR-RR-RRRRRRRRC1CRMVkOF0HMCR8OsDNNF0HMMRHR Q  0R18jR4(.n3-g4gnR
RRRRRR-R-R0hFC
#:RRRRRRRR-R-RRRRRR2RNR0)Ck#sMRR-G-R[$VRFsZRR=GRR+[R$
RLRRCMoH
RRRRRRRRR--tRC0PkNDCFRVsCRoMNCsDNRO#RC
RRRRRsRRCs0kMmRBv upX-'5Z 3),ZR-32Qv;R
RRMRC8-R""
;
RRRRVOkM0MHFR""-R:5ZRRHMBumvp_ Xuqmp)RR2skC0sBMRmpvu uX_m)pqR
H#RRRRRRRR-7-RCs#OHHb0F
M:RRRRRRRR-R-RRRRRRCR1CkRVMHO0F8MRCNODsHN0FHMRM RQ 1 R048Rj3(n.g-4gRn
RRRRR-RR-FRh0:C#
RRRRRRRRR--RRRRRNRR2CR)0Mks#ZR53tvq,3RZqR)t+qRvau]_QR2
RRRRR-RR-RRRRRRRRRL2)kC0sRM#ZMRFRsCsFRs
RRRRRPRRNNsHLRDCau v: R)q
p;RRRRLHCoMR
RRRRRR-R-RCBEOP	RN8DHHR0$FHVRM0bkRoNskMlC0R#
RRRRRHRRVRR5Z)3qtRR=-avq]Q_uR02RE
CMRRRRRRRRRRRRRRRRR#RN#0CsRpwq1R 
RRRRRRRRRRRRRRRRRRRRRRRRRsRRCsbF0ZR"3tq)R-=Rv]qa_RuQH-MR5"Z2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRP#CC0sH$)R );m)
RRRRRRRRRRRRRRRRsRRCs0kM;RZ
RRRRRRRR8CMR;HV
R
RRRRRR-R-R0tCRHbsMbOHNPDRNCDkRsVFRMoCCDsNR#ONCR
RRRRRR Rav:uR= R)q5p'Z)3qt+2RRavq]Q_u;R

RRRRRsRRCs0kMmRBv upXm_up'q)5vZ3qRt,t_ auh)QBqQupq_ep5z au v2
2;RRRRCRM8";-"
R
RRkRVMHO0FBMRmRhK5RZ:HBMRmpvu RX2skC0sBMRmpvu HXR#R
RRRRRR-R-R#7CObsH0MHF:R
RRRRRR-R-RRRRRRRR1RCCVOkM0MHFRO8CDNNs0MHFRRHMQ   R810R(4jn-3.4ngg
RRRRRRRRR--hCF0#R:
RRRRR-RR-RRRRRRRRRN2)kC0sRM#GRR-[V$RFZsRRG=RR[+R$R
RRCRLo
HMRRRRRRRR-t-RCP0RNCDkRsVFRMoCCDsNR#ONCR
RRRRRRCRs0MksRvBmuXp '35Z)R ,-QZ3v
2;RRRRCRM8BKmh;R

RVRRk0MOHRFMBKmhR:5ZRRHMBumvp_ Xuqmp)s2RCs0kMmRBv upXm_upRq)HR#
RRRRR-RR-CR7#HOsbF0HMR:
RRRRR-RR-RRRRRRRRC1CRMVkOF0HMCR8OsDNNF0HMMRHR Q  0R18jR4(.n3-g4gnR
RRRRRR-R-R0hFC
#:RRRRRRRR-R-RRRRRR2RNR0)Ck#sMRvBmuXp RMOF[Nko05CRZq3vt-,RZ)3qtR2
RRRRR-RR-RRRRRRRRRL2)kC0sRM#ZMRFRsCsFRs
RRRRR-RR-R
RRRRRRNRPsLHNDaCR :vuRQu)huBQqep_q pz;R
RRCRLo
HMRRRRRRRR-B-RE	CORDPNH08H$VRFRbHMkN0RslokC#M0
RRRRRRRRRHV53RZqR)t=vR-q_a]u2QRRC0EMR
RRRRRRRRRRRRRRRRRNC##sw0Rq p1
RRRRRRRRRRRRRRRRRRRRRRRRRRRRbsCFRs0"qZ3)=tRRq-vau]_QMRHRhBmK25Z"R
RRRRRRRRRRRRRRRRRRRRRRRRRRCR#PHCs0 $R)))m;R
RRRRRRRRRRRRRRRRRskC0sZMR;R
RRRRRRMRC8VRH;R

RRRRR-RR-CRt0sRbHHMObRNDPkNDCFRVsCRoMNCsDNRO#RC
RRRRRHRRVRR5Z)3qtRR=v]qa_RuQFZsR3tq)Rj=R32jRRC0EMR
RRRRRRRRRRRRRR Rav:uR=3RZq;)t
RRRRRRRR#CDCR
RRRRRRRRRRRRRR Rav:uR=ZR-3tq);R
RRRRRRMRC8VRH;R

RRRRRRRRskC0sBMRmpvu uX_m)pq'35Zv,qtRva u
2;RRRRCRM8BKmh;R

RVRRk0MOHRFM1aT)5RZ:HBMRmpvu 2XRR0sCkRsMBumvpR XHR#
RRRRR-RR-CR7#HOsbF0HMR:
RRRRR-RR-RRRRRRRRC1CRMVkOF0HMCR8OsDNNF0HMMRHR Q  0R18jR4(.n3-g4gnR
RRRRRR-R-R0hFC
#:RRRRRRRR-R-RRRRRRFRhMRC
RRRRRPRRNNsHLRDCZva uRR:Bumvp_ Xuqmp)R;
RRRRRPRRNNsHLRDCZamzRB:Rmpvu 
X;RRRRRRRRPHNsNCLDRqavtRR:)p q;R
RRRRRRNRPsLHNDaCRqR)t: R)q
p;RRRRLHCoMR
RRRRRR-R-R0tCRDPNkVCRF#sRbHCONODRN##C
RRRRRRRRRHV5RRZ=qRvaB]_Zm )R02RE
CMRRRRRRRRRRRRRRRRskC0svMRq_a]B)Z mR;
RRRRRCRRMH8RV
;
RRRRRRRR-t-RCP0RNCDkRsVFRMoCCDsNR#ONCR
RRRRRRaRZ Rvu:B=Rmpvu aX_mm_up5q)Z
2;RRRRRRRRatvqRR:=1aT)5 Zavvu3q;t2
RRRRRRRR)aqt=R:R6j3* Zavqu3)
t;
RRRRRRRRRHV5mRB1q5a)Rt2>3RjjRR20MEC
RRRRRRRRRRRRRRRRzZma 3)RR:=atvq*1Bm5)aqt
2;RRRRRRRRRRRRRRRRZamz3RQv:a=Rv*qt15Qhatq)2R;
RRRRRRRRRRRRRsRRCs0kMmRZz
a;RRRRRRRRCRM8H
V;
RRRRRRRRRHV5mRB1q5a)Rt2<3RjjRR20MEC
RRRRRRRRRRRRRRRRzZma 3)RR:=atvq*1Bm5)aqtRR+v]qa_2uQ;R
RRRRRRRRRRRRRRmRZzQa3v=R:RqavtQ*1hq5a)+tRRavq]Q_u2R;
RRRRRRRRRRRRRsRRCs0kMmRZz
a;RRRRRRRRCRM8H
V;
RRRRRRRRRHV5QR1hq5a)Rt2>3RjjRR20MEC
RRRRRRRRRRRRRRRRzZma 3)RR:=j;3j
RRRRRRRRRRRRRRRRzZmav3QRR:=atvq*h1Q5)aqt
2;RRRRRRRRRRRRRRRRskC0sZMRm;za
RRRRRRRR8CMR;HV
R
RRRRRRmRZz)a3 =R:Rjj3;R
RRRRRRmRZzQa3v=R:RqavtQ*1hq5a)+tRRavq]Q_u2R;
RRRRRsRRCs0kMmRZz
a;RRRRCRM81aT);R

RVRRk0MOHRFM1aT)5RZ:HBMRmpvu uX_m)pqRs2RCs0kMmRBv upXm_upRq)HR#
RRRRR-RR-CR7#HOsbF0HMR:
RRRRR-RR-RRRRRRRRC1CRMVkOF0HMCR8OsDNNF0HMMRHR Q  0R18jR4(.n3-g4gnR
RRRRRR-R-R0hFC
#:RRRRRRRR-R-RRRRRR2RNR0)Ck#sMRFZRMsRCs
Fs
RRRRRRRRsPNHDNLCmRZz:aRRvBmuXp _pumq
);RRRRRRRRPHNsNCLDRqavtRR:)p q;R
RRRRRRNRPsLHNDaCRqR)t: R)q
p;RRRRLHCoMR
RRRRRR-R-RCBEOP	RN8DHHR0$FHVRM0bkRoNskMlC0R#
RRRRRHRRVRR5Z)3qtRR=-avq]Q_uR02RE
CMRRRRRRRRRRRRRRRRR#RN#0CsRpwq1R 
RRRRRRRRRRRRRRRRRRRRRRRRRsRRCsbF0ZR"3tq)R-=Rv]qa_RuQH1MRT5)aZ
2"RRRRRRRRRRRRRRRRRRRRRRRRRRRR#CCPs$H0R) )m
);RRRRRRRRRRRRRRRRRCRs0MksR
Z;RRRRRRRRCRM8H
V;
RRRRRRRRR--tRC0PkNDCFRVsbR#CNOHDNRO#
C#RRRRRRRRH5VRRvZ3q=tRRjj3R8NMRqZ3)=tRRjj3R02RE
CMRRRRRRRRRRRRRRRRskC0sZMR;R
RRRRRRMRC8VRH;R

RRRRR-RR-CRt0sRbHHMObRNDPkNDCFRVsCRoMNCsDNRO#RC
RRRRRaRRvRqt:1=RT5)aZq3vt
2;RRRRRRRRatq)RR:=j*36Z)3qt
;
RRRRRRRRZamz3tvqRR:=uQm1a Qe_q) pa'5v2qt;R

RRRRRHRRVRR5B5m1atq)2RR<jR3j2ER0CRM
RRRRRRRRRRRRRaRRqR)t:a=RqR)t+qRvau]_QR;
RRRRRCRRMH8RV
;
RRRRRRRRH5VRRm5B1q5a)Rt2=3RjjN2RM58R15Qhatq)2RR<j23jR02RE
CMRRRRRRRRRRRRRRRRatq)RR:=atq)Rv+Rq_a]u
Q;RRRRRRRRCRM8H
V;
RRRRRRRRzZma)3qt=R:Rat _Qu)huBQqep_q pz5)aqt
2;RRRRRRRRskC0sZMRm;za
RRRR8CMR)1Ta
;
RRRRVOkM0MHFRu X5RZ:HBMRmpvu 2XRR0sCkRsMBumvpR XHR#
RRRRR-RR-CR7#HOsbF0HMR:
RRRRR-RR-RRRRRRRRC1CRMVkOF0HMCR8OsDNNF0HMMRHR Q  0R18jR4(.n3-g4gnR
RRRRRR-R-R0hFC
#:RRRRRRRR-R-RRRRRRFRhM
C
RRRRRRRRPHNsNCLDRva u):R ;qp
RRRRoLCHRM
RRRRR-RR-CRt0NRPDRkCVRFs#ObCHRNDOCN##R
RRRRRRVRHRZ5RRv=Rq_a]B)Z mRR20MEC
RRRRRRRRRRRRRRRR0sCkRsMv]qa_qBA14 _;R
RRRRRRMRC8VRH;R

RRRRRHRRVRR5Z 3)Rj=R32jRRC0EMR
RRRRRRRRRRRRRRVRHRZ5R3RQv=qRvau]_QsRFRQZ3vRR=-avq]Q_uR02RE
CMRRRRRRRRRRRRRRRRRRRRRRRRskC0sBMRmpvu 5X'-j43,3Rjj
2;RRRRRRRRRRRRRRRRCRM8H
V;
RRRRRRRRRRRRRRRRRHV53RZQ=vRRavq]Q_u_ me)R_.2ER0CRM
RRRRRRRRRRRRRRRRRRRRRsRRCs0kMqRvaB]_A q1_
K;RRRRRRRRRRRRRRRRCRM8H
V;
RRRRRRRRRRRRRRRRRHV53RZQ=vRRq-vau]_Qe_m .)_R02RE
CMRRRRRRRRRRRRRRRRRRRRRRRRskC0sBMRmpvu 5X'j,3jR3-4j
2;RRRRRRRRRRRRRRRRCRM8H
V;RRRRRRRRCRM8H
V;
RRRRRRRRR--tRC0PkNDCFRVsCRoMNCsDNRO#RC
RRRRRaRR Rvu: =RXZu532) ;R
RRRRRRCRs0MksRvBmuXp ' 5avBu*mZ1532Qv, Rav1u*QZh532Qv2R;
RCRRM 8RX
u;
RRRRMVkOF0HMXR u:5ZRRHMBumvp_ Xuqmp)RR2skC0sBMRmpvu uX_m)pqR
H#RRRRRRRR-7-RCs#OHHb0F
M:RRRRRRRR-R-RRRRRRCR1CkRVMHO0F8MRCNODsHN0FHMRM RQ 1 R048Rj3(n.g-4gRn
RRRRR-RR-FRh0:C#
RRRRRRRRR--RRRRRNRR2CR)0Mks#RRZFCMRsssF
R
RRRRRRNRPsLHNDZCRau vRB:Rmpvu 
X;RRRRRRRRPHNsNCLDRl0Cb):R ;qp
RRRRRRRRsPNHDNLCmRZz:aRRvBmuXp _pumq
);RRRRLHCoMR
RRRRRR-R-RCBEOP	RN8DHHR0$FHVRM0bkRoNskMlC0R#
RRRRRHRRVRR5Z)3qtRR=-avq]Q_uR02RE
CMRRRRRRRRRRRRRRRRR#RN#0CsRpwq1R 
RRRRRRRRRRRRRRRRRRRRRRRRRsRRCsbF0ZR"3tq)R-=Rv]qa_RuQH MRXZu52R"
RRRRRRRRRRRRRRRRRRRRRRRRR#RRCsPCHR0$ m)))R;
RRRRRRRRRRRRRRRRR0sCkRsMZR;
RRRRRCRRMH8RV
;
RRRRRRRR-t-RCP0RNCDkRsVFRC#bODHNR#ONCR#
RRRRRHRRVRR5Zq3vtRR=jR3jNRM8Z)3qtRR=jR3j2ER0CRM
RRRRRRRRRRRRRsRRCs0kMmRBv upXm_up'q)5j43,3Rjj
2;RRRRRRRRCRM8H
V;
RRRRRRRRRHV53RZvRqt=qRvau]_QMRN8ZR53tq)Rv=Rq_a]umQ_e_ ).sRF
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR3RZqR)t=vR-q_a]umQ_e_ ).2R2RC0EMR
RRRRRRRRRRRRRRCRs0MksRvBmuXp _pumq5)'4,3jRavq]Q_u2R;
RRRRRCRRMH8RV
;
RRRRRRRRH5VRRvZ3q=tRRavq]Q_u_ me)R_.2ER0CRM
RRRRRRRRRRRRRHRRVRR5Z)3qtRR=v]qa__uQm)e _2.RRC0EMR
RRRRRRRRRRRRRRRRRRRRRRCRs0MksRvBmuXp _pumq5)'4,3jRavq]Q_u_ me)2_.;R
RRRRRRRRRRRRRRMRC8VRH;R

RRRRRRRRRRRRRHRRVRR5Z)3qtRR=-avq]Q_u_ me)R_.2ER0CRM
RRRRRRRRRRRRRRRRRRRRRsRRCs0kMmRBv upXm_up'q)5j43,vR-q_a]umQ_e_ ).
2;RRRRRRRRRRRRRRRRCRM8H
V;RRRRRRRRCRM8H
V;
RRRRRRRRR--tRC0bMsHONHbDNRPDRkCVRFsoCCMsRNDOCN#
RRRRRRRR Zav:uR=mRup_q)aBm_mpvu ZX52R;
RRRRRZRRm3zavRqt:u=Rma1QQ_e )p q'X5 ua5Z 3vu)2 2;R
RRRRRRmRZzqa3):tR= Rta)_uQQhBu_qpezqp a5Z 3vuQ;v2
R
RRRRRRCRs0MksRzZmaR;
RCRRM 8RX
u;
RRRRMVkOF0HMmRpt:5ZRRHMBumvpR X2CRs0MksRvBmuXp R
H#RRRRRRRR-7-RCs#OHHb0F
M:RRRRRRRR-R-RRRRRRCR1CkRVMHO0F8MRCNODsHN0FHMRM RQ 1 R048Rj3(n.g-4gRn
RRRRR-RR-FRh0:C#
RRRRRRRRR--RRRRRNRR2CR)0Mks#mRBv upX)'5 'qpp,mWRjj32MRFRsCsF
s
RRRRRRRRPHNsNCLDR Zav:uRRvBmuXp _pumq
);RRRRRRRRPHNsNCLDRva uRR:)p q;R
RRCRLo
HMRRRRRRRR-B-RE	CORDPNH08H$VRFRbHMkN0RslokC#M0
RRRRRRRRRHV53RZ)= RRjj3RMRN83RZQ=vRRjj3R02RE
CMRRRRRRRRRRRRRRRRNC##sw0Rq p1
RRRRRRRRRRRRRRRRRRRRRRRRbsCFRs0")Z3 RR=jR3jNRM8Zv3QRj=R3HjRMmRpt25Z"R
RRRRRRRRRRRRRRRRRRRRRRCR#PHCs0 $R)))m;R
RRRRRRRRRRRRRRCRs0MksRvBmuXp ' 5)qpp'mRW,j23j;R
RRRRRRMRC8VRH;R

RRRRR-RR-CRt0NRPDRkCVRFs#ObCHRNDOCN##R
RRRRRRVRHRZ5R3RQv=3RjjRR20MEC
RRRRRRRRRRRRRRRRRHV53RZ)= RR3-4jRR20MEC
RRRRRRRRRRRRRRRRRRRRRRRR0sCkRsMBumvp' X5jj3,qRvau]_Q
2;RRRRRRRRRRRRRRRRCRM8H
V;RRRRRRRRRRRRRRRRH5VRR)Z3 RR=v]qa_2 RRC0EMR
RRRRRRRRRRRRRRRRRRRRRRCRs0MksRavq]A_Bq_1 4R;
RRRRRRRRRRRRRCRRMH8RVR;
RRRRRRRRRRRRRHRRVRR5Z 3)R4=R32jRRC0EMR
RRRRRRRRRRRRRRRRRRRRRRCRs0MksRavq]Z_B ;)m
RRRRRRRRRRRRRRRR8CMR;HV
RRRRRRRR8CMR;HV
R
RRRRRRVRHRZ5R3R) =3RjjRR20MEC
RRRRRRRRRRRRRRRRRHV5QZ3vRR=423jRC0EMR
RRRRRRRRRRRRRRRRRRRRRRCRs0MksRvBmuXp '35jjv,Rq_a]umQ_e_ ).
2;RRRRRRRRRRRRRRRRCRM8H
V;RRRRRRRRRRRRRRRRH5VRZv3QR-=R423jRC0EMR
RRRRRRRRRRRRRRRRRRRRRRCRs0MksRvBmuXp '35jj-,Rv]qa__uQm)e _;.2
RRRRRRRRRRRRRRRR8CMR;HV
RRRRRRRR8CMR;HV
R
RRRRRR-R-R0tCRDPNkVCRFosRCsMCNODRN
#CRRRRRRRRZva u=R:RvBmuXp __amuqmp)25Z;R
RRRRRR Rav:uR=mRpta5Z 3vuv2qt;R
RRRRRRCRs0MksRvBmuXp ' 5avRu,Zva u)3qt
2;RRRRCRM8p;mt
R
RRkRVMHO0FpMRm5t.ZH:RMmRBv upXRR2skC0sBMRmpvu HXR#R
RRRRRR-R-R#7CObsH0MHF:R
RRRRRR-R-RRRRRRRR1RCCVOkM0MHFRO8CDNNs0MHFRRHMQ   R810R(4jn-3.4ngg
RRRRRRRRR--hCF0#R:
RRRRR-RR-RRRRRRRRRN2)kC0sRM#Bumvp' X5q) pm'pWj,R3Rj2FCMRsssF
R
RRRRRRNRPsLHNDZCRau vRB:Rmpvu uX_m)pq;R
RRRRRRNRPsLHNDaCR Rvu: R)q
p;RRRRLHCoMR

RRRRR-RR-ERBCRO	PHND8$H0RRFVHkMb0sRNoCklM
0#RRRRRRRRH5VRR)Z3 RR=jR3jR8NMRQZ3vRR=jR3j2ER0CRM
RRRRRRRRRRRRRNRR#s#C0qRwp
1 RRRRRRRRRRRRRRRRRRRRRRRRsFCbs"0RZ 3)Rj=R3NjRMZ8R3RQv=3RjjMRHRtpm.25Z"R
RRRRRRRRRRRRRRRRRRRRRRCR#PHCs0 $R)))m;R
RRRRRRRRRRRRRRCRs0MksRvBmuXp ' 5)qpp'mRW,j23j;R
RRRRRRMRC8VRH;R

RRRRR-RR-CRt0NRPDRkCVRFs#ObCHRNDOCN##R
RRRRRRVRHRZ5R3RQv=3RjjRR20MEC
RRRRRRRRRRRRRRRRRHV53RZ)= RRj.3R02RE
CMRRRRRRRRRRRRRRRRRRRRRRRRskC0svMRq_a]B1Aq ;_4
RRRRRRRRRRRRRRRR8CMR;HV
RRRRRRRRRRRRRRRRRHV53RZ)= RRj43R02RE
CMRRRRRRRRRRRRRRRRRRRRRRRRskC0svMRq_a]B)Z mR;
RRRRRRRRRRRRRCRRMH8RVR;
RRRRRCRRMH8RV
;
RRRRRRRR-t-RCP0RNCDkRsVFRMoCCDsNR#ONCR
RRRRRRaRZ Rvu:B=Rmpvu aX_mm_up5q)Z
2;RRRRRRRRau vRR:=v]qa_tpm.w_m_p *mZt5au v3tvq2R;
RRRRRsRRCs0kMmRBv upXa'5 ,vuRavq]m_ptm._w*_ Zva u)3qt
2;RRRRCRM8p.mt;R

RVRRk0MOHRFMp4mtj:5ZRRHMBumvpR X2CRs0MksRvBmuXp R
H#RRRRRRRR-7-RCs#OHHb0F
M:RRRRRRRR-R-RRRRRRCR1CkRVMHO0F8MRCNODsHN0FHMRM RQ 1 R048Rj3(n.g-4gRn
RRRRR-RR-FRh0:C#
RRRRRRRRR--RRRRRNRR2CR)0Mks#mRBv upX)'5 'qpp,mWRjj32MRFRsCsF
s
RRRRRRRRPHNsNCLDR Zav:uRRvBmuXp _pumq
);RRRRRRRRPHNsNCLDRva uRR:)p q;R
RRCRLo
HMRRRRRRRR-B-RE	CORDPNH08H$VRFRbHMkN0RslokC#M0
RRRRRRRRRHV53RZ)= RRjj3RMRN83RZQ=vRRjj3R02RE
CMRRRRRRRRRRRRRRRRNC##sw0Rq p1
RRRRRRRRRRRRRRRRRRRRRRRRbsCFRs0")Z3 RR=jR3jNRM8Zv3QRj=R3HjRMmRpt54jZ
2"RRRRRRRRRRRRRRRRRRRRRRRR#CCPs$H0R) )m
);RRRRRRRRRRRRRRRRskC0sBMRmpvu 5X')p q'Wpm,3Rjj
2;RRRRRRRRCRM8H
V;
RRRRRRRRR--tRC0PkNDCFRVsbR#CNOHDNRO#
C#RRRRRRRRH5VRRQZ3vRR=jR3j2ER0CRM
RRRRRRRRRRRRRHRRVRR5Z 3)R4=RjR3j2ER0CRM
RRRRRRRRRRRRRRRRRRRRRsRRCs0kMqRvaB]_A q1_
4;RRRRRRRRRRRRRRRRCRM8H
V;RRRRRRRRRRRRRRRRH5VRR)Z3 RR=4R3j2ER0CRM
RRRRRRRRRRRRRRRRRRRRRsRRCs0kMqRvaB]_Zm );R
RRRRRRRRRRRRRRMRC8VRH;R
RRRRRRMRC8VRH;R

RRRRR-RR-CRt0NRPDRkCVRFsoCCMsRNDOCN#
RRRRRRRR Zav:uR=mRBv upXm_a_pumqZ)52R;
RRRRRaRR Rvu:v=Rq_a]p4mtjw_m_p *mZt5au v3tvq2R;
RRRRRsRRCs0kMmRBv upXa'5 ,vuRavq]m_pt_4jm w_* Zavqu3);t2
RRRR8CMRtpm4
j;
R
RRkRVMHO0FpMRmZt5:MRHRvBmuXp _pumq2)RR0sCkRsMBumvp_ Xuqmp)#RH
RRRRRRRRR--7OC#s0HbH:FM
RRRRRRRRR--RRRRR1RRCVCRk0MOHRFM8DCON0sNHRFMHQMR R  1R084nj(34.-g
gnRRRRRRRR-h-RF#0C:R
RRRRRR-R-RRRRRRRRN)2RCs0kMB#Rmpvu uX_m)pq5q) pQ']tR],v]qa_2uQRRFMCFsssR

RRRRRPRRNNsHLRDCZva uRR:Bumvp; X
RRRRRRRRsPNHDNLCmRZz:aRRvBmuXp _pumq
);RRRRLHCoMR
RRRRRR-R-RCBEOP	RN8DHHR0$FHVRM0bkRoNskMlC0R#
RRRRRHRRVRR5Zq3vt=R<Rjj3R02RE
CMRRRRRRRRRRRRRRRRNC##sw0Rq p1
RRRRRRRRRRRRRRRRRRRRRRRRbsCFRs0"vZ3q<tR=3RjjMRHRtpm5"Z2
RRRRRRRRRRRRRRRRRRRRRRRRP#CC0sH$)R );m)
RRRRRRRRRRRRRRRR0sCkRsMBumvp_ Xuqmp))'5 'qp]]Qt,qRvau]_Q
2;RRRRRRRRCRM8H
V;
RRRRRRRRRHV53RZqR)t=vR-q_a]u2QRRC0EMR
RRRRRRRRRRRRRRRRRNC##sw0Rq p1
RRRRRRRRRRRRRRRRRRRRRRRRRRRRbsCFRs0"qZ3)=tRRq-vau]_QMRHRtpm5"Z2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRP#CC0sH$)R );m)
RRRRRRRRRRRRRRRR0sCkRsMBumvp_ Xuqmp))'5 'qp]]Qt,qRvau]_Q
2;RRRRRRRRCRM8H
V;
RRRRRRRRR--BbFlkR0CPkNDCFRVsbR#CNOHDNRO#
C#RRRRRRRRH5VRZq3vtRR=4R3j2ER0CRM
RRRRRRRRRRRRRHRRVRR5Z)3qtRR=jR3j2ER0CRM
RRRRRRRRRRRRRRRRRRRRRsRRCs0kMmRBv upXm_up'q)5jj3,3Rjj
2;RRRRRRRRRRRRRRRRCRM8H
V;
RRRRRRRRRRRRRRRRRHV53RZqR)t=qRvau]_QRR20MEC
RRRRRRRRRRRRRRRRRRRRRRRR0sCkRsMBumvp_ Xuqmp)v'5q_a]uRQ,v]qa__uQm)e _;.2
RRRRRRRRRRRRRRRR8CMR;HV
R
RRRRRRRRRRRRRRVRHRZ5R3tq)Rv=Rq_a]umQ_e_ ).RR20MEC
RRRRRRRRRRRRRRRRRRRRRRRR0sCkRsMBumvp_ Xuqmp)v'5q_a]umQ_e_ ).v,Rq_a]umQ_e_ ).
2;RRRRRRRRRRRRRRRRCRM8H
V;
RRRRRRRRRRRRRRRRRHV53RZqR)t=vR-q_a]umQ_e_ ).RR20MEC
RRRRRRRRRRRRRRRRRRRRRRRR0sCkRsMBumvp_ Xuqmp)v'5q_a]umQ_e_ ).-,Rv]qa__uQm)e _;.2
RRRRRRRRRRRRRRRR8CMR;HV
RRRRRRRR8CMR;HV
R
RRRRRRVRHRZ5R3tvqRv=Rq_a] MRN83RZqR)t=3RjjRR20MEC
RRRRRRRRRRRRRRRR0sCkRsMBumvp_ Xuqmp)4'53Rj,j23j;R
RRRRRRMRC8VRH;R

RRRRR-RR-FRBl0bkCNRPDRkCVRFsoCCMsRNDOCN#
RRRRRRRR Zav)u3 =R:Rtpm5vZ3q;t2
RRRRRRRR ZavQu3v=R:RqZ3)
t;RRRRRRRRZamzRR:=Bumvp_ Xaum_m)pq5 Zav;u2
RRRRRRRR0sCkRsMZamz;R
RRMRC8mRpt
;

R
RRkRVMHO0FpMRm5t.ZH:RMmRBv upXm_upRq)2CRs0MksRvBmuXp _pumqH)R#R
RRRRRR-R-R#7CObsH0MHF:R
RRRRRR-R-RRRRRRRR1RCCVOkM0MHFRO8CDNNs0MHFRRHMQ   R810R(4jn-3.4ngg
RRRRRRRRR--hCF0#R:
RRRRR-RR-RRRRRRRRRN2)kC0sRM#Bumvp_ Xuqmp) 5)q]p'Q,t]Ravq]Q_u2MRFRsCsF
s
RRRRRRRRPHNsNCLDR Zav:uRRvBmuXp ;R
RRRRRRNRPsLHNDZCRmRza:mRBv upXm_up;q)
RRRRoLCHRM
RRRRR-RR-ERBCRO	PHND8$H0RRFVHkMb0sRNoCklM
0#RRRRRRRRH5VRRvZ3q<tR=3RjjRR20MEC
RRRRRRRRRRRRRRRR#N#CRs0w1qp R
RRRRRRRRRRRRRRRRRRRRRRCRsb0FsR3"ZvRqt<j=R3HjRMmRptZ.52R"
RRRRRRRRRRRRRRRRRRRRR#RRCsPCHR0$ m)))R;
RRRRRRRRRRRRRsRRCs0kMmRBv upXm_up'q)5q) pQ']tR],v]qa_2uQ;R
RRRRRRMRC8VRH;R

RRRRRHRRVRR5Z)3qtRR=-avq]Q_uR02RE
CMRRRRRRRRRRRRRRRRR#RN#0CsRpwq1R 
RRRRRRRRRRRRRRRRRRRRRRRRRsRRCsbF0ZR"3tq)R-=Rv]qa_RuQHpMRm5t.Z
2"RRRRRRRRRRRRRRRRRRRRRRRRRRRR#CCPs$H0R) )m
);RRRRRRRRRRRRRRRRskC0sBMRmpvu uX_m)pq' 5)q]p'Q,t]Ravq]Q_u2R;
RRRRRCRRMH8RV
;
RRRRRRRR-B-RFklb0PCRNCDkRsVFRC#bODHNR#ONCR#
RRRRRHRRVZR53tvqR4=R3NjRMZ8R3tq)Rj=R32jRRC0EMR
RRRRRRRRRRRRRRCRs0MksRvBmuXp _pumq5)'j,3jRjj32R;
RRRRRCRRMH8RV
;
RRRRRRRRH5VRRvZ3q=tRRj.3R8NMRqZ3)=tRRjj3R02RE
CMRRRRRRRRRRRRRRRRskC0sBMRmpvu uX_m)pq'354jj,R3;j2
RRRRRRRR8CMR;HV
R
RRRRRR-R-RlBFbCk0RDPNkVCRFosRCsMCNODRN
#CRRRRRRRRZva u 3)RR:=v]qa_tpm.w_m_p *mZt53tvq2R;
RRRRRZRRau v3RQv:v=Rq_a]p.mt__mw 3*Zq;)t
RRRRRRRRzZma=R:RvBmuXp __amuqmp)a5Z 2vu;R
RRRRRRCRs0MksRzZmaR;
RCRRMp8Rm;t.
R
RRkRVMHO0FpMRmjt45RZ:HBMRmpvu uX_m)pqRs2RCs0kMmRBv upXm_upRq)HR#
RRRRR-RR-CR7#HOsbF0HMR:
RRRRR-RR-RRRRRRRRC1CRMVkOF0HMCR8OsDNNF0HMMRHR Q  0R18jR4(.n3-g4gnR
RRRRRR-R-R0hFC
#:RRRRRRRR-R-RRRRRR2RNR0)Ck#sMRvBmuXp _pumq))5 'qp]]Qt,qRvau]_QF2RMsRCs
FsRRRRRRRRPHNsNCLDR Zav:uRRvBmuXp ;R
RRRRRRNRPsLHNDZCRmRza:mRBv upXm_up;q)
RRRRoLCHRM
RRRRR-RR-ERBCRO	PHND8$H0RRFVHkMb0sRNoCklM
0#RRRRRRRRH5VRRvZ3q<tR=3RjjRR20MEC
RRRRRRRRRRRRRRRR#N#CRs0w1qp R
RRRRRRRRRRRRRRRRRRRRRRCRsb0FsR3"ZvRqt<j=R3HjRMmRpt54jZ
2"RRRRRRRRRRRRRRRRRRRRRRRR#CCPs$H0R) )m
);RRRRRRRRRRRRRRRRskC0sBMRmpvu uX_m)pq' 5)q]p'Q,t]Ravq]Q_u2R;
RRRRRCRRMH8RV
;

RRRRRRRRRHV53RZqR)t=vR-q_a]u2QRRC0EMR
RRRRRRRRRRRRRRRRRNC##sw0Rq p1
RRRRRRRRRRRRRRRRRRRRRRRRRRRsFCbs"0RZ)3qtRR=-avq]Q_uRRHMp4mtj25Z"R
RRRRRRRRRRRRRRRRRRRRRRRRRRP#CC0sH$)R );m)
RRRRRRRRRRRRRRRR0sCkRsMBumvp_ Xuqmp))'5 'qp]]Qt,qRvau]_Q
2;RRRRRRRRCRM8H
V;
RRRRRRRRR--BbFlkR0CPkNDCFRVsbR#CNOHDNRO#
C#RRRRRRRRH5VRZq3vtRR=4R3jNRM8Z)3qtRR=jR3j2ER0CRM
RRRRRRRRRRRRRsRRCs0kMmRBv upXm_up'q)5jj3,3Rjj
2;RRRRRRRRCRM8H
V;
RRRRRRRRRHV53RZvRqt=jR43NjRMZ8R3tq)Rj=R32jRRC0EMR
RRRRRRRRRRRRRRCRs0MksRvBmuXp _pumq5)'4,3jRjj32R;
RRRRRCRRMH8RV
;
RRRRRRRR-B-RFklb0PCRNCDkRsVFRMoCCDsNR#ONCR
RRRRRRaRZ 3vu): R=qRvap]_mjt4__mw m*pt35Zv2qt;R
RRRRRRaRZ 3vuQ:vR=qRvap]_mjt4__mw 3*Zq;)t
RRRRRRRRzZma=R:RvBmuXp __amuqmp)a5Z 2vu;R
RRRRRRCRs0MksRzZmaR;
RCRRMp8Rmjt4;R

RVRRk0MOHRFMp5mtZH:RMmRBv upXA;Rq:1 RRHM)p qRs2RCs0kMmRBv upX#RH
RRRRRRRRR--7OC#s0HbH:FM
RRRRRRRRR--RRRRR1RRCVCRk0MOHRFM8DCON0sNHRFMHQMR R  1R084nj(34.-g
gnRRRRRRRR-h-RF#0C:R
RRRRRR-R-RRRRRRRRN)2RCs0kMB#Rmpvu 5X')p q'Wpm,3RjjF2RMsRCs
Fs
RRRRRRRRsPNHDNLCaRZ Rvu:mRBv upXm_up;q)
RRRRRRRRsPNHDNLC Rav u)R):R ;qp
RRRRRRRRsPNHDNLC RavvuQR):R ;qp
RRRRoLCHRM
RRRRR-RR-ERBCRO	PHND8$H0RRFVHkMb0sRNoCklM
0#RRRRRRRRH5VRR)Z3 RR=jR3jR8NMRQZ3vRR=jR3j2ER0CRM
RRRRRRRRRRRRRNRR#s#C0qRwp
1 RRRRRRRRRRRRRRRRRRRRRRRRsFCbs"0RZ 3)Rj=R3NjRMZ8R3RQv=3RjjMRHRtpm5AZ,q21 "R
RRRRRRRRRRRRRRRRRRRRRRCR#PHCs0 $R)))m;R
RRRRRRRRRRRRRRCRs0MksRvBmuXp ' 5)qpp'mRW,j23j;R
RRRRRRMRC8VRH;R

RRRRRHRRVRR5A q1RR<=jR3jFAsRqR1 =3R4jRR20MEC
RRRRRRRRRRRRRRRR#N#CRs0w1qp R
RRRRRRRRRRRRRRRRRRRRRRCRsb0FsRq"A1< R=3RjjsRFR1Aq RR=4R3jHpMRmZt5,1Aq 
2"RRRRRRRRRRRRRRRRRRRRRRRR#CCPs$H0R) )m
);RRRRRRRRRRRRRRRRskC0sBMRmpvu 5X')p q'Wpm,3Rjj
2;RRRRRRRRCRM8H
V;
RRRRRRRRR--tRC0PkNDCFRVsbR#CNOHDNRO#
C#RRRRRRRRH5VRRQZ3vRR=jR3j2ER0CRM
RRRRRRRRRRRRRHRRVRR5Z 3)RA=RqR1 2ER0CRM
RRRRRRRRRRRRRRRRRRRRRsRRCs0kMqRvaB]_A q1_
4;RRRRRRRRRRRRRRRRCRM8H
V;RRRRRRRRRRRRRRRRH5VRR)Z3 RR=4R3j2ER0CRM
RRRRRRRRRRRRRRRRRRRRRsRRCs0kMqRvaB]_Zm );R
RRRRRRRRRRRRRRMRC8VRH;R
RRRRRRMRC8VRH;R

RRRRR-RR-CRt0NRPDRkCVRFsoCCMsRNDOCN#
RRRRRRRR Zav:uR=mRBv upXm_a_pumqZ)52R;
RRRRRaRR )vu =R:Rtpm5 Zavvu3qRt,A q12R;
RRRRRaRR Qvuv=R:R Zavqu3)pt/mAt5q21 ;R
RRRRRRCRs0MksRvBmuXp ' 5av u), RavvuQ2R;
RCRRMp8Rm
t;
RRRRMVkOF0HMmRpt:5ZRRHMBumvp_ Xuqmp)A;Rq:1 RRHM)p qRs2RCs0kMmRBv upXm_upRq)HR#
RRRRR-RR-CR7#HOsbF0HMR:
RRRRR-RR-RRRRRRRRC1CRMVkOF0HMCR8OsDNNF0HMMRHR Q  0R18jR4(.n3-g4gnR
RRRRRR-R-R0hFC
#:RRRRRRRR-R-RRRRRR2RNR0)Ck#sMRvBmuXp _pumq))5 'qp]]Qt,qRvau]_QF2RMsRCs
Fs
RRRRRRRRsPNHDNLCaRZ Rvu:mRBv upXR;
RRRRRPRRNNsHLRDCZamzRB:Rmpvu uX_m)pq;R
RRCRLo
HMRRRRRRRR-B-RE	CORDPNH08H$VRFRbHMkN0RslokC#M0
RRRRRRRRRHV53RZvRqt<j=R32jRRC0EMR
RRRRRRRRRRRRRR#RN#0CsRpwq1R 
RRRRRRRRRRRRRRRRRRRRRsRRCsbF0ZR"3tvqRR<=jR3jHpMRmZt5,1Aq 
2"RRRRRRRRRRRRRRRRRRRRRRRR#CCPs$H0R) )m
);RRRRRRRRRRRRRRRRskC0sBMRmpvu uX_m)pq' 5)q]p'Q,t]Ravq]Q_u2R;
RRRRRCRRMH8RV
;
RRRRRRRRH5VRR1Aq =R<Rjj3RRFsA q1R4=R32jRRC0EMR
RRRRRRRRRRRRRR#RN#0CsRpwq1R 
RRRRRRRRRRRRRRRRRRRRRsRRCsbF0AR"qR1 <j=R3FjRsqRA1= RRj43RRHMp5mtZq,A1" 2
RRRRRRRRRRRRRRRRRRRRRRRRP#CC0sH$)R );m)
RRRRRRRRRRRRRRRR0sCkRsMBumvp_ Xuqmp))'5 'qp]]Qt,qRvau]_Q
2;RRRRRRRRCRM8H
V;
RRRRRRRRRHV53RZqR)t=vR-q_a]u2QRRC0EMR
RRRRRRRRRRRRRR#RN#0CsRpwq1R 
RRRRRRRRRRRRRRRRRRRRRRRRRCRsb0FsR3"ZqR)t=vR-q_a]uHQRMmRpt,5ZA q12R"
RRRRRRRRRRRRRRRRRRRRRRRRRCR#PHCs0 $R)))m;R
RRRRRRRRRRRRRRCRs0MksRvBmuXp _pumq5)')p q't]Q]v,Rq_a]u;Q2
RRRRRRRR8CMR;HV
R
RRRRRR-R-RlBFbCk0RDPNkVCRF#sRbHCONODRN##C
RRRRRRRRRHV5vZ3q=tRRj43R8NMRqZ3)=tRRjj3R02RE
CMRRRRRRRRRRRRRRRRskC0sBMRmpvu uX_m)pq'35jjj,R3;j2
RRRRRRRR8CMR;HV
R
RRRRRRVRHRZ5R3tvqRA=RqR1 NRM8Z)3qtRR=jR3j2ER0CRM
RRRRRRRRRRRRRsRRCs0kMmRBv upXm_up'q)5j43,3Rjj
2;RRRRRRRRCRM8H
V;
RRRRRRRRR--BbFlkR0CPkNDCFRVsCRoMNCsDNRO#RC
RRRRRZRRau v3R) :p=RmZt53tvq,qRA1; 2
RRRRRRRR ZavQu3v=R:RqZ3)pt/mAt5q21 ;R
RRRRRRmRZz:aR=mRBv upXm_a_pumqZ)5au v2R;
RRRRRsRRCs0kMmRZz
a;RRRRCRM8p;mt
R

RVRRk0MOHRFM15QhZH:RMmRBv upXRR2skC0sBMRmpvu HXR#R
RRRRRR-R-R#7CObsH0MHF:R
RRRRRR-R-RRRRRRRR1RCCVOkM0MHFRO8CDNNs0MHFRRHMQ   R810R(4jn-3.4ngg
RRRRRRRRR--hCF0#R:
RRRRR-RR-RRRRRRRRMhFCR
RRCRLo
HMRRRRRRRR-t-RCP0RNCDkRsVFRC#bODHNR#ONCR#
RRRRRHRRVRR5Zv3QRj=R32jRRC0EMR
RRRRRRRRRRRRRRVRHRZ5R3R) =3RjjsRFR)Z3 RR=v]qa_2uQRC0EMR
RRRRRRRRRRRRRRRRRRRRRRCRs0MksRavq]Z_B ;)m
RRRRRRRRRRRRRRRR8CMR;HV
RRRRRRRR8CMR;HV
R
RRRRRR-R-R0tCRDPNkVCRFosRCsMCNODRN
#CRRRRRRRRskC0sBMRmpvu 5X'15QhZ 3)2m*B1Z]532Qv,mRB135Z)* 21]Qh5QZ3v;22
RRRR8CMRh1Q;R

RVRRk0MOHRFM15QhZH:RMmRBv upXm_upRq)2CRs0MksRvBmuXp _pumqH)R#R
RRRRRR-R-R#7CObsH0MHF:R
RRRRRR-R-RRRRRRRR1RCCVOkM0MHFRO8CDNNs0MHFRRHMQ   R810R(4jn-3.4ngg
RRRRRRRRR--hCF0#R:
RRRRR-RR-RRRRRRRRRN2)kC0sRM#Bumvp_ Xuqmp)35jjj,R3Rj2FCMRsssF
R
RRRRRRNRPsLHNDZCR4Z,R.RR:Bumvp; X
RRRRRRRRsPNHDNLCmRZz:aRRvBmuXp _pumq
);RRRRLHCoMR
RRRRRR-R-RCBEOP	RN8DHHR0$FHVRM0bkRoNskMlC0R#
RRRRRHRRVRR5Z)3qtRR=-avq]Q_uR02RE
CMRRRRRRRRRRRRRRRRNC##sw0Rq p1
RRRRRRRRRRRRRRRRRRRRRRRRRRRRbsCFRs0"qZ3)=tRRq-vau]_QMRHRh1Q5"Z2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRP#CC0sH$)R );m)
RRRRRRRRRRRRRRRR0sCkRsMBumvp_ Xuqmp)j'53Rj,j23j;R
RRRRRRMRC8VRH;R

RRRRR-RR-FRBl0bkCNRPDRkCVRFs#ObCHRNDOCN##R
RRRRRRVRHRZ5R3tvqRj=R3NjRMZ8R3tq)Rj=R32jRRC0EMR
RRRRRRRRRRRRRRCRs0MksRvBmuXp _pumq5)'j,3jRjj32R;
RRRRRCRRMH8RV
;
RRRRRRRRH5VRRvZ3q=tRRavq]Q_uR8NMRqZ3)=tRRjj3R02RE
CMRRRRRRRRRRRRRRRRskC0sBMRmpvu uX_m)pq'35jjj,R3;j2
RRRRRRRR8CMR;HV
R
RRRRRR-R-RlBFbCk0RDPNkVCRFosRCsMCNODRN
#CRRRRRRRRZ:4R=mRup_q)aBm_mpvu ZX52R;
RRRRRZRR.=R:RvBmuXp 'Q51h45Z32) *1Bm]45Z32Qv,mRB145Z32) *h1Q]45Z32Qv2R;
RRRRRZRRmRza:B=Rmpvu aX_mm_up5q)Z;.2
RRRRRRRR0sCkRsMZamz;R
RRMRC8QR1h
;
RRRRVOkM0MHFR1Bm5RZ:HBMRmpvu 2XRR0sCkRsMBumvpR XHR#
RRRRR-RR-CR7#HOsbF0HMR:
RRRRR-RR-RRRRRRRRC1CRMVkOF0HMCR8OsDNNF0HMMRHR Q  0R18jR4(.n3-g4gnR
RRRRRR-R-R0hFC
#:RRRRRRRR-R-RRRRRRFRhMRC
RLRRCMoH
R

RRRRR-RR-CRt0NRPDRkCVRFs#ObCHRNDOCN##R
RRRRRRVRHRZ5R3RQv=3RjjRR20MEC
RRRRRRRRRRRRRRRRRHV53RZ)= RRavq]Q_u_ me)R_.FZsR3R) =vR-q_a]umQ_e_ ).02RE
CMRRRRRRRRRRRRRRRRRRRRRRRRskC0svMRq_a]B)Z mR;
RRRRRRRRRRRRRCRRMH8RVR;
RRRRRCRRMH8RV
;
RRRRRRRR-t-RCP0RNCDkRsVFRMoCCDsNR#ONCR
RRRRRRCRs0MksRvBmuXp 'm5B135Z)* 2B]m15QZ3vR2,-h1Q5)Z3 12*Q5h]Zv3Q2
2;RRRRCRM8B;m1
R
RRkRVMHO0FBMRmZ15:MRHRvBmuXp _pumq2)RR0sCkRsMBumvp_ Xuqmp)#RH
RRRRRRRRR--7OC#s0HbH:FM
RRRRRRRRR--RRRRR1RRCVCRk0MOHRFM8DCON0sNHRFMHQMR R  1R084nj(34.-g
gnRRRRRRRR-h-RF#0C:R
RRRRRR-R-RRRRRRRRN)2RCs0kMB#Rmpvu uX_m)pq5jj3,3RjjF2RMsRCs
Fs
RRRRRRRRsPNHDNLC4RZ,.RZRB:Rmpvu 
X;RRRRRRRRPHNsNCLDRzZmaRR:Bumvp_ Xuqmp)R;
RLRRCMoH
RRRRRRRRR--BOEC	NRPDHH80F$RVMRHbRk0Nksol0CM#R
RRRRRRVRHRZ5R3tq)R-=Rv]qa_RuQ2ER0CRM
RRRRRRRRRRRRRNRR#s#C0qRwp
1 RRRRRRRRRRRRRRRRRRRRRRRRRRRRsFCbs"0RZ)3qtRR=-avq]Q_uRRHMB5m1Z
2"RRRRRRRRRRRRRRRRRRRRRRRRRRRR#CCPs$H0R) )m
);RRRRRRRRRRRRRRRRskC0sBMRmpvu uX_m)pq'35jjj,R3;j2
RRRRRRRR8CMR;HV
R
RRRRRR-R-RlBFbCk0RDPNkVCRF#sRbHCONODRN##C
RRRRRRRRRHV53RZvRqt=qRvau]_Qe_m .)_R8NMRqZ3)=tRRjj3R02RE
CMRRRRRRRRRRRRRRRRskC0sBMRmpvu uX_m)pq'35jjj,R3;j2
RRRRRRRR8CMR;HV
R
RRRRRRVRHRZ5R3tvqRv=Rq_a]umQ_e_ ).MRN83RZqR)t=qRvau]_QRR20MEC
RRRRRRRRRRRRRRRR0sCkRsMBumvp_ Xuqmp)j'53Rj,j23j;R
RRRRRRMRC8VRH;R

RRRRR-RR-FRBl0bkCNRPDRkCVRFsoCCMsRNDOCN#
RRRRRRRRRZ4:u=Rm)pq__amBumvp5 XZ
2;RRRRRRRRZ:.R=mRBv upXB'5mZ154 3)2m*B1Z]54v3Q2-,R15QhZ)43 12*Q5h]ZQ43v;22
RRRRRRRRzZma=R:RvBmuXp __amuqmp).5Z2R;
RRRRRsRRCs0kMmRZz
a;RRRRCRM8B;m1
R
RRkRVMHO0F1MRQ5h]ZH:RMmRBv upXRR2skC0sBMRmpvu HXR#R
RRRRRR-R-R#7CObsH0MHF:R
RRRRRR-R-RRRRRRRR1RCCVOkM0MHFRO8CDNNs0MHFRRHMQ   R810R(4jn-3.4ngg
RRRRRRRRR--hCF0#R:
RRRRR-RR-RRRRRRRRMhFCR
RRCRLo
HMRRRRRRRR-t-RCP0RNCDkRsVFRC#bODHNR#ONCR#
RRRRRHRRVRR5Z 3)Rj=R32jRRC0EMR
RRRRRRRRRRRRRRVRHRZ5R3RQv=3RjjsRFRQZ3vRR=v]qa_RuQ2ER0CRM
RRRRRRRRRRRRRRRRRRRRRsRRCs0kMqRvaB]_Zm );R
RRRRRRRRRRRRRRMRC8VRH;



RRRRRRRRRRRRRRRRRHV53RZQ=vRRavq]Q_u_ me)R_.2ER0CRM
RRRRRRRRRRRRRRRRRRRRRsRRCs0kMqRvaB]_A q1_
K;RRRRRRRRRRRRRRRRCRM8H
V;
RRRRRRRRRRRRRRRRRHV53RZQ=vRRq-vau]_Qe_m .)_R02RE
CMRRRRRRRRRRRRRRRRRRRRRRRRskC0s-MRv]qa_qBA1K _;R
RRRRRRRRRRRRRRMRC8VRH;R
RRRRRRMRC8VRH;R

RRRRR-RR-CRt0NRPDRkCVRFsoCCMsRNDOCN#
RRRRRRRR0sCkRsMBumvp' X5h1Q]35Z)* 2B5m1Zv3Q2B,Rm51]Z 3)2Q*1h35ZQ2v2;R
RRMRC8QR1h
];
RRRRMVkOF0HMQR1hZ]5:MRHRvBmuXp _pumq2)RR0sCkRsMBumvp_ Xuqmp)#RH
RRRRRRRRR--7OC#s0HbH:FM
RRRRRRRRR--RRRRR1RRCVCRk0MOHRFM8DCON0sNHRFMHQMR R  1R084nj(34.-g
gnRRRRRRRR-h-RF#0C:R
RRRRRR-R-RRRRRRRRN)2RCs0kMB#Rmpvu uX_m)pq5jj3,3RjjF2RMsRCs
Fs
RRRRRRRRsPNHDNLC4RZ,.RZRB:Rmpvu 
X;RRRRRRRRPHNsNCLDRzZmaRR:Bumvp_ Xuqmp)R;
RLRRCMoH
RRRRRRRRR--BOEC	NRPDHH80F$RVMRHbRk0Nksol0CM#R
RRRRRRVRHRZ5R3tq)R-=Rv]qa_RuQ2ER0CRM
RRRRRRRRRRRRRNRR#s#C0qRwp
1 RRRRRRRRRRRRRRRRRRRRRRRRRRRRsFCbs"0RZ)3qtRR=-avq]Q_uRRHM1]Qh5"Z2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRP#CC0sH$)R );m)
RRRRRRRRRRRRRRRR0sCkRsMBumvp_ Xuqmp)j'53Rj,j23j;R
RRRRRRMRC8VRH;R

RRRRR-RR-FRBl0bkCNRPDRkCVRFs#ObCHRNDOCN##R
RRRRRRVRHRZ5R3tvqRj=R3NjRMZ8R3tq)Rj=R32jRRC0EMR
RRRRRRRRRRRRRRCRs0MksRvBmuXp _pumq5)'j,3jRjj32R;
RRRRRCRRMH8RV
;
RRRRRRRRH5VRRvZ3q=tRRavq]Q_uR8NMRqZ3)=tRRavq]Q_u_ me)R_.2ER0CRM
RRRRRRRRRRRRRsRRCs0kMmRBv upXm_up'q)5jj3,3Rjj
2;RRRRRRRRCRM8H
V;
RRRRRRRRRHV53RZvRqt=qRvau]_Qe_m .)_R8NMRqZ3)=tRRavq]Q_u_ me)R_.2ER0CRM
RRRRRRRRRRRRRsRRCs0kMmRBv upXm_up'q)5j43,qRvau]_Qe_m .)_2R;
RRRRRCRRMH8RV
;
RRRRRRRRH5VRRvZ3q=tRRavq]Q_u_ me)R_.NRM8Z)3qtRR=-avq]Q_u_ me)R_.2ER0CRM
RRRRRRRRRRRRRsRRCs0kMmRBv upXm_up'q)5j43,vR-q_a]umQ_e_ ).
2;RRRRRRRRCRM8H
V;
RRRRRRRRR--BbFlkR0CPkNDCFRVsCRoMNCsDNRO#RC
RRRRRZRR4=R:Rpumqa)_mm_Bv upX25Z;R
RRRRRR.RZRR:=Bumvp' X5h1Q]45Z32) *1Bm53Z4Q,v2R1Bm]45Z32) *h1Q53Z4Q2v2;R
RRRRRRmRZz:aR=mRBv upXm_a_pumqZ)5.
2;RRRRRRRRskC0sZMRm;za
RRRR8CMRh1Q]
;

RRRRMVkOF0HMmRB1Z]5:MRHRvBmuXp Rs2RCs0kMmRBv upX#RH
RRRRRRRRR--7OC#s0HbH:FM
RRRRRRRRR--RRRRR1RRCVCRk0MOHRFM8DCON0sNHRFMHQMR R  1R084nj(34.-g
gnRRRRRRRR-h-RF#0C:R
RRRRRR-R-RRRRRRRRhCFM
RRRRoLCHRM
RRRRR-RR-CRt0NRPDRkCVRFs#ObCHRNDOCN##R
RRRRRRVRHRZ5R3R) =3RjjRR20MEC
RRRRRRRRRRRRRRRRRHV53RZQ=vRRjj3R02RE
CMRRRRRRRRRRRRRRRRRRRRRRRRskC0svMRq_a]B1Aq ;_4
RRRRRRRRRRRRRRRR8CMR;HV
R
RRRRRRRRRRRRRRVRHRZ5R3RQv=qRvau]_QRR20MEC
RRRRRRRRRRRRRRRRRRRRRRRR0sCkRsM-avq]A_Bq_1 4R;
RRRRRRRRRRRRRCRRMH8RV
;
RRRRRRRRRRRRRRRRH5VRRQZ3vRR=v]qa__uQm)e _F.Rs3RZQ=vRRq-vau]_Qe_m .)_R02RE
CMRRRRRRRRRRRRRRRRRRRRRRRRskC0svMRq_a]B)Z mR;
RRRRRRRRRRRRRCRRMH8RVR;
RRRRRCRRMH8RV
;
RRRRRRRR-t-RCP0RNCDkRsVFRMoCCDsNR#ONCR
RRRRRRCRs0MksRvBmuXp 'm5B1Z]532) *1Bm5QZ3vR2,1]Qh5)Z3 12*QZh532Qv2R;
RCRRMB8Rm;1]
R
RRkRVMHO0FBMRm51]ZH:RMmRBv upXm_upRq)2CRs0MksRvBmuXp _pumqH)R#R
RRRRRR-R-R#7CObsH0MHF:R
RRRRRR-R-RRRRRRRR1RCCVOkM0MHFRO8CDNNs0MHFRRHMQ   R810R(4jn-3.4ngg
RRRRRRRRR--hCF0#R:
RRRRR-RR-RRRRRRRRRN2)kC0sRM#Bumvp_ Xuqmp)35jjj,R3Rj2FCMRsssF
R
RRRRRRNRPsLHNDZCR4Z,R.RR:Bumvp; X
RRRRRRRRsPNHDNLCmRZz:aRRvBmuXp _pumq
);RRRRLHCoMR
RRRRRR-R-RCBEOP	RN8DHHR0$FHVRM0bkRoNskMlC0R#
RRRRRHRRVRR5Z)3qtRR=-avq]Q_uR02RE
CMRRRRRRRRRRRRRRRRNC##sw0Rq p1
RRRRRRRRRRRRRRRRRRRRRRRRRRRRbsCFRs0"qZ3)=tRRq-vau]_QMRHR1Bm]25Z"R
RRRRRRRRRRRRRRRRRRRRRRRRRRCR#PHCs0 $R)))m;R
RRRRRRRRRRRRRRCRs0MksRvBmuXp _pumq5)'j,3jRjj32R;
RRRRRCRRMH8RV
;
RRRRRRRR-B-RFklb0PCRNCDkRsVFRC#bODHNR#ONCR#
RRRRRHRRVRR5Zq3vtRR=jR3jNRM8Z)3qtRR=jR3j2ER0CRM
RRRRRRRRRRRRRsRRCs0kMmRBv upXm_up'q)5j43,3Rjj
2;RRRRRRRRCRM8H
V;
RRRRRRRRRHV53RZvRqt=qRvau]_QMRN83RZqR)t=qRvau]_Qe_m .)_R02RE
CMRRRRRRRRRRRRRRRRskC0sBMRmpvu uX_m)pq'354jv,Rq_a]u;Q2
RRRRRRRR8CMR;HV
R
RRRRRRVRHRZ5R3tvqRv=Rq_a]umQ_e_ ).MRN83RZqR)t=qRvau]_Qe_m .)_R02RE
CMRRRRRRRRRRRRRRRRskC0sBMRmpvu uX_m)pq'35jjj,R3;j2
RRRRRRRR8CMR;HV
R
RRRRRRVRHRZ5R3tvqRv=Rq_a]umQ_e_ ).MRN83RZqR)t=vR-q_a]umQ_e_ ).RR20MEC
RRRRRRRRRRRRRRRR0sCkRsMBumvp_ Xuqmp)j'53Rj,j23j;R
RRRRRRMRC8VRH;R

RRRRR-RR-FRBl0bkCNRPDRkCVRFsoCCMsRNDOCN#
RRRRRRRRRZ4:u=Rm)pq__amBumvp5 XZ
2;RRRRRRRRZ:.R=mRBv upXB'5m51]Z)43 B2*mZ154v3Q21,RQ5h]Z)43 12*QZh54v3Q2
2;RRRRRRRRZamzRR:=Bumvp_ Xaum_m)pq52Z.;R
RRRRRRCRs0MksRzZmaR;
RCRRMB8Rm;1]
R

R-RR-R
RR-R-RHqs0CEl0RHOmsbCNs0F#R
RR-R-
RRRRMVkOF0HM+R""RR5pH:RMmRBv upXR;R)H:RMmRBv upXRR2skC0sBMRmpvu HXR#R
RRRRRR-R-R#7CObsH0MHF:R
RRRRRR-R-RRRRRRRR1RCCVOkM0MHFRO8CDNNs0MHFRRHMQ   R810R(4jn-3.4ngg
RRRRRRRRR--hCF0#R:
RRRRR-RR-RRRRRRRRMhFCR
RRCRLo
HMRRRRRRRRskC0sBMRmpvu 5X'p 3)R)+R3,) RQp3vRR+)v3Q2R;
RCRRM"8R+
";
RRRRMVkOF0HM+R""RR5pH:RM R)qRp;)H:RMmRBv upXRR2skC0sBMRmpvu HXR#R
RRRRRR-R-R#7CObsH0MHF:R
RRRRRR-R-RRRRRRRR1RCCVOkM0MHFRO8CDNNs0MHFRRHMQ   R810R(4jn-3.4ngg
RRRRRRRRR--hCF0#R:
RRRRR-RR-RRRRRRRRMhFCR
RRCRLo
HMRRRRRRRRskC0sBMRmpvu 5X'pRR+) 3),3R)Q;v2
RRRR8CMR""+;R

RVRRk0MOHRFM"R+"5:RpRRHMBumvp; XR:R)RRHM)p qRR2RRCRs0MksRvBmuXp R
H#RRRRRRRR-7-RCs#OHHb0F
M:RRRRRRRR-R-RRRRRRCR1CkRVMHO0F8MRCNODsHN0FHMRM RQ 1 R048Rj3(n.g-4gRn
RRRRR-RR-FRh0:C#
RRRRRRRRR--RRRRRhRRF
MCRRRRLHCoMR
RRRRRRCRs0MksRvBmuXp '35p)+ RRR),pv3Q2R;
RCRRM"8R+
";
RRRRMVkOF0HM+R""pR5:MRHRvBmuXp _pumqR);)H:RMmRBv upXm_up2q)
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR0sCkRsMBumvp_ Xuqmp)#RH
RRRRRRRRR--7OC#s0HbH:FM
RRRRRRRRR--RRRRR1RRCVCRk0MOHRFM8DCON0sNHRFMHQMR R  1R084nj(34.-g
gnRRRRRRRR-h-RF#0C:R
RRRRRR-R-RRRRRRRRN)2RCs0kMB#Rmpvu uX_m)pq'35jjj,R3Rj2FCMRsssF
RRRRRRRR
--RRRRRRRRPHNsNCLDR,ZpRRZ):mRBv upXR;
RRRRRPRRNNsHLRDCZamzRB:Rmpvu uX_m)pq;R
RRCRLo
HMRRRRRRRR-B-RE	CORDPNH08H$VRFRbHMkN0RslokC#M0
RRRRRRRRRHV53RpqR)t=vR-q_a]u2QRRC0EMR
RRRRRRRRRRRRRR#RN#0CsRpwq1R 
RRRRRRRRRRRRRRRRRRRRRRRRRsRRCsbF0pR"3tq)R-=Rv]qa_RuQH+MR5)p,2R"
RRRRRRRRRRRRRRRRRRRRRRRRR#RRCsPCHR0$ m)))R;
RRRRRRRRRRRRRsRRCs0kMmRBv upXm_up'q)5jj3,3Rjj
2;RRRRRRRRCRM8H
V;
R
RRRRRRVRHR)5R3tq)R-=Rv]qa_RuQ2ER0CRM
RRRRRRRRRRRRRNRR#s#C0qRwp
1 RRRRRRRRRRRRRRRRRRRRRRRRRRRRsFCbs"0R))3qtRR=-avq]Q_uRRHM+,5p)
2"RRRRRRRRRRRRRRRRRRRRRRRRRRRR#CCPs$H0R) )m
);RRRRRRRRRRRRRRRRskC0sBMRmpvu uX_m)pq'35jjj,R3;j2
RRRRRRRR8CMR;HV
R
RRRRRR-R-R0tCRHbsMbOHNPDRNCDk
RRRRRRRRRZp:u=Rm)pq__amBumvp5 XR2pR;R
RRRRRR)RZRR:=uqmp)m_a_vBmuXp 5RR)2R;
RRRRRZRRmRza:B=Rmpvu aX_mm_up5q)Bumvp' X53Zp)+ RR3Z))R ,ZQp3vZR+)v3Q2
2;RRRRRRRRskC0sZMRm;za
RRRR8CMR""+;R

RVRRk0MOHRFM"R+"5:RpRRHM)p q;)RR:MRHRvBmuXp _pumqR)2skC0sBMRmpvu uX_m)pqR
H#RRRRRRRR-7-RCs#OHHb0F
M:RRRRRRRR-R-RRRRRRCR1CkRVMHO0F8MRCNODsHN0FHMRM RQ 1 R048Rj3(n.g-4gRn
RRRRR-RR-FRh0:C#
RRRRRRRRR--RRRRRNRR2CR)0Mks#mRBv upXm_up'q)5jj3,3RjjF2RMsRCs
FsRRRRRRRRPHNsNCLDRRZ):mRBv upXR;
RRRRRPRRNNsHLRDCZamzRB:Rmpvu uX_m)pq;R
RRCRLo
HMRRRRRRRR-B-RE	CORDPNH08H$VRFRbHMkN0RslokC#M0
RRRRRRRRRHV53R)qR)t=vR-q_a]u2QRRC0EMR
RRRRRRRRRRRRRR#RN#0CsRpwq1R 
RRRRRRRRRRRRRRRRRRRRRRRRRsRRCsbF0)R"3tq)R-=Rv]qa_RuQH+MR5)p,2R"
RRRRRRRRRRRRRRRRRRRRRRRRR#RRCsPCHR0$ m)))R;
RRRRRRRRRRRRRsRRCs0kMmRBv upXm_up'q)5jj3,3Rjj
2;RRRRRRRRCRM8H
V;
RRRRRRRRR--tRC0bMsHONHbDNRPD
kCRRRRRRRRZ:)R=mRup_q)aBm_mpvu RX5);R2
RRRRRRRRzZma=R:RvBmuXp __amuqmp)m5Bv upXp'5RZ+R) 3),)RZ32Qv2R;
RRRRRsRRCs0kMmRZz
a;RRRRCRM8";+"
R
RRkRVMHO0F"MR+5"RRRp:HBMRmpvu uX_m)pq;)RR:MRHRq) ps2RCs0kMmRBv upXm_upRq)HR#
RRRRR-RR-CR7#HOsbF0HMR:
RRRRR-RR-RRRRRRRRC1CRMVkOF0HMCR8OsDNNF0HMMRHR Q  0R18jR4(.n3-g4gnR
RRRRRR-R-R0hFC
#:RRRRRRRR-R-RRRRRR2RNR0)Ck#sMRvBmuXp _pumq5)'j,3jRjj32MRFRsCsFRs
RRRRR-RR-R
RRRRRRNRPsLHNDZCRpRR:Bumvp; X
RRRRRRRRsPNHDNLCmRZz:aRRvBmuXp _pumq
);RRRRLHCoMR
RRRRRR-R-RCBEOP	RN8DHHR0$FHVRM0bkRoNskMlC0R#
RRRRRHRRVRR5p)3qtRR=-avq]Q_uR02RE
CMRRRRRRRRRRRRRRRRNC##sw0Rq p1
RRRRRRRRRRRRRRRRRRRRRRRRRRRRbsCFRs0"qp3)=tRRq-vau]_QMRHRp+5,")2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRP#CC0sH$)R );m)
RRRRRRRRRRRRRRRR0sCkRsMBumvp_ Xuqmp)j'53Rj,j23j;R
RRRRRRMRC8VRH;R

RRRRR-RR-CRt0sRbHHMObRNDPkNDCR
RRRRRRpRZRR:=uqmp)m_a_vBmuXp 5RRp2R;
RRRRRZRRmRza:B=Rmpvu aX_mm_up5q)Bumvp' X53Zp)+ RRR),ZQp3v;22
RRRRRRRR0sCkRsMZamz;R
RRMRC8+R""
;
RRRRVOkM0MHFR""-Rp5R:MRHRvBmuXp ;)RR:MRHRvBmuXp Rs2RCs0kMmRBv upX#RH
RRRRRRRRR--7OC#s0HbH:FM
RRRRRRRRR--RRRRR1RRCVCRk0MOHRFM8DCON0sNHRFMHQMR R  1R084nj(34.-g
gnRRRRRRRR-h-RF#0C:R
RRRRRR-R-RRRRRRRRhCFM
RRRRoLCHRM
RRRRRsRRCs0kMmRBv upXp'53R) -3R))R ,pv3QR)-R32Qv;R
RRMRC8-R""
;
RRRRVOkM0MHFR""-Rp5R:MRHRq) pR;RR)RR:MRHRvBmuXp Rs2RCs0kMmRBv upX#RH
RRRRRRRRR--7OC#s0HbH:FM
RRRRRRRRR--RRRRR1RRCVCRk0MOHRFM8DCON0sNHRFMHQMR R  1R084nj(34.-g
gnRRRRRRRR-h-RF#0C:R
RRRRRR-R-RRRRRRRRhCFM
RRRRoLCHRM
RRRRRsRRCs0kMmRBv upXp'5R)-R3,) R3-4jRR*)v3Q2R;
RCRRM"8R-
";
RRRRMVkOF0HM-R""RR5pH:RMmRBv upXR;R)H:RM R)q2pRRRRRskC0sBMRmpvu HXR#R
RRRRRR-R-R#7CObsH0MHF:R
RRRRRR-R-RRRRRRRR1RCCVOkM0MHFRO8CDNNs0MHFRRHMQ   R810R(4jn-3.4ngg
RRRRRRRRR--hCF0#R:
RRRRR-RR-RRRRRRRRMhFCR
RRCRLo
HMRRRRRRRRskC0sBMRmpvu 5X'p 3)R)-R,3RpQ;v2
RRRR8CMR""-;R

RVRRk0MOHRFM"R-"5:RpRRHMBumvp_ Xuqmp));R:MRHRvBmuXp _pumq
)2RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRskC0sBMRmpvu uX_m)pqR
H#RRRRRRRR-7-RCs#OHHb0F
M:RRRRRRRR-R-RRRRRRCR1CkRVMHO0F8MRCNODsHN0FHMRM RQ 1 R048Rj3(n.g-4gRn
RRRRR-RR-FRh0:C#
RRRRRRRRR--RRRRRNRR2CR)0Mks#mRBv upXm_up'q)5jj3,3RjjF2RMsRCs
FsRRRRRRRR-R-
RRRRRPRRNNsHLRDCZRp,Z:)RRvBmuXp ;R
RRRRRRNRPsLHNDZCRmRza:mRBv upXm_up;q)
RRRRoLCHRM
RRRRR-RR-ERBCRO	PHND8$H0RRFVHkMb0sRNoCklM
0#RRRRRRRRH5VRRqp3)=tRRq-vau]_QRR20MEC
RRRRRRRRRRRRRRRR#N#CRs0w1qp R
RRRRRRRRRRRRRRRRRRRRRRRRRRCRsb0FsR3"pqR)t=vR-q_a]uHQRM5R-p2,)"R
RRRRRRRRRRRRRRRRRRRRRRRRRRCR#PHCs0 $R)))m;R
RRRRRRRRRRRRRRCRs0MksRvBmuXp _pumq5)'j,3jRjj32R;
RRRRRCRRMH8RV
;
RRRRRRRRH5VRRq)3)=tRRq-vau]_QRR20MEC
RRRRRRRRRRRRRRRR#N#CRs0w1qp R
RRRRRRRRRRRRRRRRRRRRRRRRRRCRsb0FsR3")qR)t=vR-q_a]uHQRM5R-p2,)"R
RRRRRRRRRRRRRRRRRRRRRRRRRRCR#PHCs0 $R)))m;R
RRRRRRRRRRRRRRCRs0MksRvBmuXp _pumq5)'j,3jRjj32R;
RRRRRCRRMH8RVR;
RRRRR-RR-CRt0sRbHHMObRNDPkNDCR
RRRRRRpRZRR:=uqmp)m_a_vBmuXp 5RRp2R;
RRRRRZRR)=R:Rpumqa)_mm_Bv upX)5RR
2;RRRRRRRRZamzRR:=Bumvp_ Xaum_m)pq5vBmuXp 'p5Z3R) -)RZ3,) R3ZpQ-vRZQ)3v;22
RRRRRRRR0sCkRsMZamz;R
RRMRC8-R""
;
RRRRVOkM0MHFR""-Rp5R:MRHRq) pR;R)H:RMmRBv upXm_up2q)R0sCkRsMBumvp_ Xuqmp)#RH
RRRRRRRRR--7OC#s0HbH:FM
RRRRRRRRR--RRRRR1RRCVCRk0MOHRFM8DCON0sNHRFMHQMR R  1R084nj(34.-g
gnRRRRRRRR-h-RF#0C:R
RRRRRR-R-RRRRRRRRN)2RCs0kMB#Rmpvu uX_m)pq'35jjj,R3Rj2FCMRsssF
RRRRRRRR
--RRRRRRRRPHNsNCLDRRZ):mRBv upXR;
RRRRRPRRNNsHLRDCZamzRB:Rmpvu uX_m)pq;R
RRCRLo
HMRRRRRRRR-B-RE	CORDPNH08H$VRFRbHMkN0RslokC#M0
RRRRRRRRRHV53R)qR)t=vR-q_a]u2QRRC0EMR
RRRRRRRRRRRRRR#RN#0CsRpwq1R 
RRRRRRRRRRRRRRRRRRRRRRRRRsRRCsbF0)R"3tq)R-=Rv]qa_RuQH-MR5)p,2R"
RRRRRRRRRRRRRRRRRRRRRRRRR#RRCsPCHR0$ m)))R;
RRRRRRRRRRRRRsRRCs0kMmRBv upXm_up'q)5jj3,3Rjj
2;RRRRRRRRCRM8H
V;
RRRRRRRRR--tRC0bMsHONHbDNRPD
kCRRRRRRRRZ:)R=mRup_q)aBm_mpvu RX5);R2
RRRRRRRRzZma=R:RvBmuXp __amuqmp)m5Bv upXp'5RZ-R) 3),4R-3Zj*)v3Q2
2;RRRRRRRRskC0sZMRm;za
RRRR8CMR""-;R

RVRRk0MOHRFM"R-"5:RpRRHMBumvp_ Xuqmp)R;R)H:RM R)qRp2skC0sBMRmpvu uX_m)pqR
H#RRRRRRRR-7-RCs#OHHb0F
M:RRRRRRRR-R-RRRRRRCR1CkRVMHO0F8MRCNODsHN0FHMRM RQ 1 R048Rj3(n.g-4gRn
RRRRR-RR-FRh0:C#
RRRRRRRRR--RRRRRNRR2CR)0Mks#mRBv upXm_up'q)5jj3,3RjjF2RMsRCs
FsRRRRRRRR-R-
RRRRRPRRNNsHLRDCZ:pRRvBmuXp ;R
RRRRRRNRPsLHNDZCRmRza:mRBv upXm_up;q)
RRRRoLCHRM
RRRRR-RR-ERBCRO	PHND8$H0RRFVHkMb0sRNoCklM
0#RRRRRRRRH5VRRqp3)=tRRq-vau]_QRR20MEC
RRRRRRRRRRRRRRRR#N#CRs0w1qp R
RRRRRRRRRRRRRRRRRRRRRRRRRRCRsb0FsR3"pqR)t=vR-q_a]uHQRM5R-p2,)"R
RRRRRRRRRRRRRRRRRRRRRRRRRRCR#PHCs0 $R)))m;R
RRRRRRRRRRRRRRCRs0MksRvBmuXp _pumq5)'j,3jRjj32R;
RRRRRCRRMH8RV
;
RRRRRRRR-t-RCb0RsOHMHDbNRDPNkRC
RRRRRZRRp=R:Rpumqa)_mm_Bv upXp5RR
2;RRRRRRRRZamzRR:=Bumvp_ Xaum_m)pq5vBmuXp 'p5Z3R) -,R)R3ZpQ2v2;R
RRRRRRCRs0MksRzZmaR;
RCRRM"8R-
";
R
RRkRVMHO0F"MR*5"RRRp:HBMRmpvu RX;RR):HBMRmpvu 2XRR0sCkRsMBumvpR XHR#
RRRRR-RR-CR7#HOsbF0HMR:
RRRRR-RR-RRRRRRRRC1CRMVkOF0HMCR8OsDNNF0HMMRHR Q  0R18jR4(.n3-g4gnR
RRRRRR-R-R0hFC
#:RRRRRRRR-R-RRRRRRFRhMRC
RLRRCMoH
RRRRRRRR0sCkRsMBumvp' X5)p3 RR*) 3)Rp-R3RQv*3R)QRv,p 3)R)*R3RQv+3RpQ*vRR))3 
2;RRRRCRM8";*"
R

RVRRk0MOHRFM"R*"5:RpRRHM)p q;)RR:MRHRvBmuXp Rs2RCs0kMmRBv upX#RH
RRRRRRRRR--7OC#s0HbH:FM
RRRRRRRRR--RRRRR1RRCVCRk0MOHRFM8DCON0sNHRFMHQMR R  1R084nj(34.-g
gnRRRRRRRR-h-RF#0C:R
RRRRRR-R-RRRRRRRRhCFM
RRRRoLCHRM
RRRRRsRRCs0kMmRBv upXp'5R)*R3,) R*pRRQ)3v
2;RRRRCRM8";*"
R
RRkRVMHO0F"MR*5"RRRp:HBMRmpvu RX;RR):H)MR Rqp2RRRR0sCkRsMBumvpR XHR#
RRRRR-RR-CR7#HOsbF0HMR:
RRRRR-RR-RRRRRRRRC1CRMVkOF0HMCR8OsDNNF0HMMRHR Q  0R18jR4(.n3-g4gnR
RRRRRR-R-R0hFC
#:RRRRRRRR-R-RRRRRRFRhMRC
RLRRCMoH
RRRRRRRR0sCkRsMBumvp' X5)p3 RR*)p,R3RQv*2R);R
RRMRC8*R""
;
RRRRVOkM0MHFR""*Rp5R:MRHRvBmuXp _pumqR);)H:RMmRBv upXm_up2q)
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR0sCkRsMBumvp_ Xuqmp)#RH
RRRRRRRRR--7OC#s0HbH:FM
RRRRRRRRR--RRRRR1RRCVCRk0MOHRFM8DCON0sNHRFMHQMR R  1R084nj(34.-g
gnRRRRRRRR-h-RF#0C:R
RRRRRR-R-RRRRRRRRN)2RCs0kMB#Rmpvu uX_m)pq'35jjj,R3Rj2FCMRsssF
RRRRRRRR
--RRRRRRRRPHNsNCLDRzZmaRR:Bumvp_ Xuqmp)R;
RLRRCMoH
RRRRRRRRR--BOEC	NRPDHH80F$RVMRHbRk0Nksol0CM#R
RRRRRRVRHRp5R3tq)R-=Rv]qa_RuQ2ER0CRM
RRRRRRRRRRRRRNRR#s#C0qRwp
1 RRRRRRRRRRRRRRRRRRRRRRRRRRRRsFCbs"0Rp)3qtRR=-avq]Q_uRRHM*,5p)
2"RRRRRRRRRRRRRRRRRRRRRRRRRRRR#CCPs$H0R) )m
);RRRRRRRRRRRRRRRRskC0sBMRmpvu uX_m)pq'35jjj,R3;j2
RRRRRRRR8CMR;HV
R
RRRRRRVRHR)5R3tq)R-=Rv]qa_RuQ2ER0CRM
RRRRRRRRRRRRRNRR#s#C0qRwp
1 RRRRRRRRRRRRRRRRRRRRRRRRRRRRsFCbs"0R))3qtRR=-avq]Q_uRRHM*,5p)
2"RRRRRRRRRRRRRRRRRRRRRRRRRRRR#CCPs$H0R) )m
);RRRRRRRRRRRRRRRRskC0sBMRmpvu uX_m)pq'35jjj,R3;j2
RRRRRRRR8CMR;HV
R
RRRRRR-R-R0tCRHbsMbOHNPDRNCDk
RRRRRRRRzZmaq3vt=R:Rvp3q*tRRv)3q
t;RRRRRRRRZamz3tq)RR:=t_ auh)QBqQupq_ep5z p)3qtRR+))3qt
2;
RRRRRRRR0sCkRsMZamz;R
RRMRC8*R""
;
RRRRVOkM0MHFR""*Rp5R:MRHRq) pR;R)H:RMmRBv upXm_up2q)R0sCkRsMBumvp_ Xuqmp)#RH
RRRRRRRRR--7OC#s0HbH:FM
RRRRRRRRR--RRRRR1RRCVCRk0MOHRFM8DCON0sNHRFMHQMR R  1R084nj(34.-g
gnRRRRRRRR-h-RF#0C:R
RRRRRR-R-RRRRRRRRN)2RCs0kMB#Rmpvu uX_m)pq'35jjj,R3Rj2FCMRsssF
RRRRRRRR
--RRRRRRRRRRRRPHNsNCLDRRZp:mRBv upXm_up;q)
RRRRRRRRsPNHDNLCmRZz:aRRvBmuXp _pumq
);RRRRLHCoMR
RRRRRR-R-RCBEOP	RN8DHHR0$FHVRM0bkRoNskMlC0R#
RRRRRHRRVRR5))3qtRR=-avq]Q_uR02RE
CMRRRRRRRRRRRRRRRRNC##sw0Rq p1
RRRRRRRRRRRRRRRRRRRRRRRRRRRRbsCFRs0"q)3)=tRRq-vau]_QMRHRp*5,")2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRP#CC0sH$)R );m)
RRRRRRRRRRRRRRRR0sCkRsMBumvp_ Xuqmp)j'53Rj,j23j;R
RRRRRRMRC8VRH;R

RRRRR-RR-CRt0sRbHHMObRNDPkNDCR
RRRRRRpRZ3tvqRR:=uQm1a Qe_q) pq'5Ap152
2;RRRRRRRRH5VRR<pRRjj3R02RE
CMRRRRRRRRRRRRRRRRZqp3):tR=qRvau]_QR;
RRRRRCRRD
#CRRRRRRRRRRRRRRRRZqp3):tR=3RjjR;
RRRRRCRRMH8RV
;
RRRRRRRRZamz3tvqRR:=Zvp3q*tRRv)3q
t;RRRRRRRRZamz3tq)RR:=t_ auh)QBqQupq_ep5z Zqp3)+tRRq)3);t2
R
RRRRRRCRs0MksRzZmaR;
RCRRM"8R*
";
RRRRMVkOF0HM*R""RR5pH:RMmRBv upXm_up;q)R:R)RRHM)p q2CRs0MksRvBmuXp _pumqH)R#R
RRRRRR-R-R#7CObsH0MHF:R
RRRRRR-R-RRRRRRRR1RCCVOkM0MHFRO8CDNNs0MHFRRHMQ   R810R(4jn-3.4ngg
RRRRRRRRR--hCF0#R:
RRRRR-RR-RRRRRRRRRN2)kC0sRM#Bumvp_ Xuqmp)j'53Rj,j23jRRFMCFsssR
RRRRRR-R-
RRRRRRRRsPNHDNLC)RZRB:Rmpvu uX_m)pq;R
RRRRRRNRPsLHNDZCRmRza:mRBv upXm_up;q)
RRRRoLCHRM
RRRRR-RR-ERBCRO	PHND8$H0RRFVHkMb0sRNoCklM
0#RRRRRRRRH5VRRqp3)=tRRq-vau]_QRR20MEC
RRRRRRRRRRRRRRRR#N#CRs0w1qp R
RRRRRRRRRRRRRRRRRRRRRRRRRRCRsb0FsR3"pqR)t=vR-q_a]uHQRM5R*p2,)"R
RRRRRRRRRRRRRRRRRRRRRRRRRRCR#PHCs0 $R)))m;R
RRRRRRRRRRRRRRCRs0MksRvBmuXp _pumq5)'j,3jRjj32R;
RRRRRCRRMH8RV
;
RRRRRRRR-t-RCb0RsOHMHDbNRDPNkRC
RRRRRZRR)q3vt=R:R1umQeaQ  _)q5p'q5A1);22
RRRRRRRRRHV5RR)<3RjjRR20MEC
RRRRRRRRRRRRRRRR3Z)qR)t:v=Rq_a]u
Q;RRRRRRRRCCD#
RRRRRRRRRRRRRRRR3Z)qR)t:j=R3
j;RRRRRRRRCRM8H
V;
RRRRRRRRzZmaq3vt=R:Rvp3q*tRR3Z)v;qt
RRRRRRRRzZma)3qt=R:Rat _Qu)huBQqep_q pz5qp3)+tRR3Z)q2)t;R

RRRRRsRRCs0kMmRZz
a;RRRRCRM8";*"
R
RRMVkOF0HM/R""RR5pH:RMmRBv upXR;R)H:RMmRBv upXRR2skC0sBMRmpvu HXR#R
RRRRRR-R-R#7CObsH0MHF:R
RRRRRR-R-RRRRRRRR1RCCVOkM0MHFRO8CDNNs0MHFRRHMQ   R810R(4jn-3.4ngg
RRRRRRRRR--hCF0#R:
RRRRR-RR-RRRRRRRRRN2)kC0sRM#Bumvp' X5q) pQ']tR],j23jRRFMCFsssR
RRRRRR-R-
RRRRRRRRsPNHDNLC Rav:uRRq) p=R:R))3 3*))+ RRQ)3v3*)Q
v;RLRRCMoH
RRRRRRRRR--BOEC	NRPDHH80F$RVMRHbRk0Nksol0CM#R
RRRRRRVRHR 5av=uRRjj32ER0CRM
RRRRRRRRRRRRRRRRNC##sw0Rq p1
RRRRRRRRRRRRRRRRRRRRRRRRbsCFRs0"0q0C0lbRR0F8HHP8BCRmpvu LXR$jR53Rj,j23j"R
RRRRRRRRRRRRRRRRRRRRRRCR#PHCs0 $R)))m;R
RRRRRRRRRRRRRRsRRCs0kMmRBv upX)'5 'qp]]Qt,3Rjj
2;RRRRRRRRCRM8H
V;
RRRRRRRRR--tRC0PkNDCR
RRRRRRCRs0MksRvBmuXp '55Rp 3)R)*R3R) +3RpQ*vRRQ)3v/2RRva uR,
RRRRRRRRRRRRRRRRRRRRRRRR5Qp3vRR*) 3)Rp-R3R) *3R)QRv2/ Rav;u2
RRRR8CMR""/;R

RkRVMHO0F"MR/5"RRRp:H)MR ;qpR:R)RRHMBumvpR X2CRs0MksRvBmuXp R
H#RRRRRRRR-7-RCs#OHHb0F
M:RRRRRRRR-R-RRRRRRCR1CkRVMHO0F8MRCNODsHN0FHMRM RQ 1 R048Rj3(n.g-4gRn
RRRRR-RR-FRh0:C#
RRRRRRRRR--RRRRRNRR2CR)0Mks#mRBv upX)'5 'qp]]Qt,3RjjF2RMsRCs
FsRRRRRRRR-R-
RRRRRPRRNNsHLRDCau vR):R Rqp:)=R3*) ) 3)R)+R3*Qv)v3Q;R
RRCRLo
HMRRRRRRRR-B-RE	CORDPNH08H$VRFRbHMkN0RslokC#M0
RRRRRRRRRHV5va uRR=j23jRC0EMR
RRRRRRRRRRRRRRNRR#s#C0qRwp
1 RRRRRRRRRRRRRRRRRRRRRRRRsFCbs"0RqC00lRb008FRH8PHCmRBv upX$RLR35jjj,R3"j2
RRRRRRRRRRRRRRRRRRRRRRRRP#CC0sH$)R );m)
RRRRRRRRRRRRRRRRCRs0MksRvBmuXp ' 5)q]p'Q,t]Rjj32R;
RRRRRCRRMH8RV
;
RRRRRRRR-t-RCP0RNCDk
RRRRRRRRva u=R:R/pRRva uR;
RRRRRsRRCs0kMBRRmpvu 5X'Rva uRR*) 3),aR- Rvu*3R)Q2vR;R
RRMRC8/R""
;
RRRRVOkM0MHFR""/Rp5R:MRHRvBmuXp ;)RR:MRHRq) pRR2RsRRCs0kMmRBv upX#RH
RRRRRRRRR--7OC#s0HbH:FM
RRRRRRRRR--RRRRR1RRCVCRk0MOHRFM8DCON0sNHRFMHQMR R  1R084nj(34.-g
gnRRRRRRRR-h-RF#0C:R
RRRRRR-R-RRRRRRRRN)2RCs0kMB#Rmpvu 5X')p q't]Q]j,R3Rj2FCMRsssF
RRRRoLCHRM
RRRRR-RR-ERBCRO	PHND8$H0RRFVHkMb0sRNoCklM
0#RRRRRRRRH5VR)RR=j23jRC0EMR
RRRRRRRRRRRRRRNRR#s#C0qRwp
1 RRRRRRRRRRRRRRRRRRRRRRRRsFCbs"0RqC00lRb008FRH8PHCmRBv upX$RLRjj3"R
RRRRRRRRRRRRRRRRRRRRRRCR#PHCs0 $R)))m;R
RRRRRRRRRRRRRRsRRCs0kMmRBv upX)'5 'qp]]Qt,3Rjj
2;RRRRRRRRCRM8H
V;
RRRRRRRRR--tRC0PkNDCR
RRRRRRCRs0MksRvBmuXp '35p)/ RRR),pv3QR)/R2R;
RCRRM"8R/
";
R
RRkRVMHO0F"MR/5"RRRp:HBMRmpvu uX_m)pq;:R)RRHMBumvp_ Xuqmp)R2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRsRRCs0kMmRBv upXm_upRq)HR#
RRRRR-RR-CR7#HOsbF0HMR:
RRRRR-RR-RRRRRRRRC1CRMVkOF0HMCR8OsDNNF0HMMRHR Q  0R18jR4(.n3-g4gnR
RRRRRR-R-R0hFC
#:RRRRRRRR-R-RRRRRR2RNR0)Ck#sMRvBmuXp _pumq5)')p q't]Q]j,R3Rj2FCMRsssF
RRRRRRRR
--RRRRRRRRPHNsNCLDRzZmaRR:Bumvp_ Xuqmp)R;
RLRRCMoH
RRRRRRRRR--BOEC	NRPDHH80F$RVMRHbRk0Nksol0CM#R
RRRRRRVRHR35)vRqt=3Rjj02RE
CMRRRRRRRRRRRRRRRRNC##sw0Rq p1
RRRRRRRRRRRRRRRRRRRRRRRRbsCFRs0"0q0C0lbRR0F8HHP8BCRmpvu uX_m)pqRRL$5jj3,3Rjj
2"RRRRRRRRRRRRRRRRRRRRRRRR#CCPs$H0R) )m
);RRRRRRRRRRRRRRRRskC0sBMRmpvu uX_m)pq' 5)q]p'Q,t]Rjj32R;
RRRRRCRRMH8RV
;
RRRRRRRRH5VRRqp3)=tRRq-vau]_QRR20MEC
RRRRRRRRRRRRRRRR#N#CRs0w1qp R
RRRRRRRRRRRRRRRRRRRRRRCRsb0FsR3"pqR)t=vR-q_a]uHQRM5R/p2,)"R
RRRRRRRRRRRRRRRRRRRRRRCR#PHCs0 $R)))m;R
RRRRRRRRRRRRRRCRs0MksRvBmuXp _pumq5)')p q't]Q]j,R3;j2
RRRRRRRR8CMR;HV
R
RRRRRRVRHR)5R3tq)R-=Rv]qa_RuQ2ER0CRM
RRRRRRRRRRRRRNRR#s#C0qRwp
1 RRRRRRRRRRRRRRRRRRRRRRRRsFCbs"0R))3qtRR=-avq]Q_uRRHM/,5p)
2"RRRRRRRRRRRRRRRRRRRRRRRR#CCPs$H0R) )m
);RRRRRRRRRRRRRRRRskC0sBMRmpvu uX_m)pq'35jjj,R3;j2
RRRRRRRR8CMR;HV
R
RRRRRR-R-R0tCRHbsMbOHNPDRNCDk
RRRRRRRRzZmaq3vt=R:Rvp3q)t/3tvq;R
RRRRRRmRZzqa3):tR= Rta)_uQQhBu_qpezqp 35pqR)t-3R)q2)t;R

RRRRRsRRCs0kMmRZz
a;RRRRCRM8";/"
R
RRkRVMHO0F"MR/5"RRRp:HBMRmpvu uX_m)pq;)RR:MRHRq) ps2RCs0kMmRBv upXm_upRq)HR#
RRRRR-RR-CR7#HOsbF0HMR:
RRRRR-RR-RRRRRRRRC1CRMVkOF0HMCR8OsDNNF0HMMRHR Q  0R18jR4(.n3-g4gnR
RRRRRR-R-R0hFC
#:RRRRRRRR-R-RRRRRR2RNR0)Ck#sMRvBmuXp _pumq5)')p q't]Q]j,R3Rj2FCMRsssF
RRRRRRRR
--RRRRRRRRPHNsNCLDRRZ):mRBv upXm_up;q)
RRRRRRRRsPNHDNLCmRZz:aRRvBmuXp _pumq
);RRRRLHCoMR
RRRRRR-R-RCBEOP	RN8DHHR0$FHVRM0bkRoNskMlC0R#
RRRRRHRRV)R5Rj=R3Rj20MEC
RRRRRRRRRRRRRRRR#N#CRs0w1qp R
RRRRRRRRRRRRRRRRRRRRRRCRsb0FsR0"q0bCl0FR0RP8HHR8CBumvp_ Xuqmp)$RLRjj3"R
RRRRRRRRRRRRRRRRRRRRRRCR#PHCs0 $R)))m;R
RRRRRRRRRRRRRRCRs0MksRvBmuXp _pumq5)')p q't]Q]j,R3;j2
RRRRRRRR8CMR;HV
R
RRRRRRVRHRp5R3tq)R-=Rv]qa_RuQ2ER0CRM
RRRRRRRRRRRRRNRR#s#C0qRwp
1 RRRRRRRRRRRRRRRRRRRRRRRRsFCbs"0Rp)3qtRR=-avq]Q_uRRHM/,5p)
2"RRRRRRRRRRRRRRRRRRRRRRRR#CCPs$H0R) )m
);RRRRRRRRRRRRRRRRskC0sBMRmpvu uX_m)pq' 5)q]p'Q,t]Rjj32R;
RRRRRCRRMH8RV
;
RRRRRRRR-t-RCb0RsOHMHDbNRDPNkRC
RRRRRZRR)q3vt=R:R1umQeaQ  _)q5p'q5A1);22
RRRRRRRRRHV)RR<jR3j0MEC
RRRRRRRRRRRRRRRR3Z)qR)t:v=Rq_a]u
Q;RRRRRRRRCCD#
RRRRRRRRRRRRRRRR3Z)qR)t:j=R3
j;RRRRRRRRCRM8H
V;
RRRRRRRRzZmaq3vt=R:Rvp3qZt/)q3vtR;
RRRRRZRRm3zaqR)t:t=R ua_)BQhQpuq_peqzp 53tq)RZ-R))3qt
2;
RRRRRRRR0sCkRsMZamz;R
RRMRC8/R""
;
RRRRVOkM0MHFR""/Rp5R:MRHRq) pR;R)H:RMmRBv upXm_up2q)R0sCkRsMBumvp_ Xuqmp)#RH
RRRRRRRRR--7OC#s0HbH:FM
RRRRRRRRR--RRRRR1RRCVCRk0MOHRFM8DCON0sNHRFMHQMR R  1R084nj(34.-g
gnRRRRRRRR-h-RF#0C:R
RRRRRR-R-RRRRRRRRN)2RCs0kMB#Rmpvu uX_m)pq' 5)q]p'Q,t]Rjj32MRFRsCsFRs
RRRRR-RR-R
RRRRRRNRPsLHNDZCRpRR:Bumvp_ Xuqmp)R;
RRRRRPRRNNsHLRDCZamzRB:Rmpvu uX_m)pq;R
RRCRLo
HMRRRRRRRR-B-RE	CORDPNH08H$VRFRbHMkN0RslokC#M0
RRRRRRRRRHV5v)3q=tRRjj32ER0CRM
RRRRRRRRRRRRRNRR#s#C0qRwp
1 RRRRRRRRRRRRRRRRRRRRRRRRsFCbs"0RqC00lRb008FRH8PHCmRBv upXm_upRq)L5$Rj,3jRjj32R"
RRRRRRRRRRRRRRRRRRRRR#RRCsPCHR0$ m)))R;
RRRRRRRRRRRRRsRRCs0kMmRBv upXm_up'q)5q) pQ']tR],j23j;R
RRRRRRMRC8VRH;R

RRRRRHRRVRR5))3qtRR=-avq]Q_uR02RE
CMRRRRRRRRRRRRRRRRNC##sw0Rq p1
RRRRRRRRRRRRRRRRRRRRRRRRbsCFRs0"q)3)=tRRq-vau]_RRHM/,5p)
2"RRRRRRRRRRRRRRRRRRRRRRRR#CCPs$H0R) )m
);RRRRRRRRRRRRRRRRskC0sBMRmpvu uX_m)pq'35jjj,R3;j2
RRRRRRRR8CMR;HV
R
RRRRRR-R-R0tCRHbsMbOHNPDRNCDk
RRRRRRRR3ZpvRqt:u=Rma1QQ_e )p q'A5q125p2R;
RRRRRHRRVRRp<3RjjER0CRM
RRRRRRRRRRRRRZRRp)3qt=R:Ravq]Q_u;R
RRRRRRDRC#RC
RRRRRRRRRRRRRZRRp)3qt=R:Rjj3;R
RRRRRRMRC8VRH;R

RRRRRZRRm3zavRqt:Z=Rpq3vt3/)v;qt
RRRRRRRRzZma)3qt=R:Rat _Qu)huBQqep_q pz53ZpqR)t-3R)q2)t;R

RRRRRsRRCs0kMmRZz
a;RRRRCRM8";/"
M
C8vRRq_a]Bumvp; X
