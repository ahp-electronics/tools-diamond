--$Header: //synplicity/map202003lat/designware/dware.vhd#1 $
@E---------------------------------------------------------------------------------------------------

---w-RHRDCRRRRR:RRRN8IsPC3E-8
-CR7#MHoRRRRRRR:B0FMN#HMRR.ULHN#OCR7#MHoWCNsRlOFbCFMMR0#
R--BbFlNRM$RRRR:$R1MHbDO$H0ROQM3-
-R07NCRRRRRRRRq:Rk.oR6.,Rj
jU-q-RkF0EsRRRR:RRRD1CPRNl)-
-RseC#MHFRRRRRd:R3-4
--
--------------------------------------------------------------------------------------------------D

HNLssQ$R ,  7)Wq k;
#QCR 3  #_08DHFoO4_4nNc3D
D;kR#C7)Wq I38_kVFM08NH_FMObFl3DND;C

M00H$WR7__VbN#88kHLR#o

CsMCH5OR
o#H_8IH0:ERR1umQeaQ =R:R;.d
bCG_8IH0:ERR1umQeaQ =R:R
U;HCCC_lOFbNDHMROC:hRQa  t)=R:R2j
;b

FRs05R
N:MRHR8#0_oDFHPO_CFO0sH5#oH_I8R0E+GRCbH_I8R0E8MFI0jFR2L;
RH:RM0R#8F_Do_HOP0COF#s5HIo_HE80RC+RGIb_HE80RI8FMR0Fj
2;sRM8:MRHR8#0_oDFHPO_CFO0sR5.8MFI0jFR2F;
bRR:H#MR0D8_FOoH;:
xR0FkR8#0_oDFHPO_CFO0sH5#oH_I8R0E+GRCbH_I8R0E8MFI0jFR2#;
0kN0#RR:FRk0#_08DHFoOC_POs0F58(RF0IMF2Rj

2;
-
-R0N0skHL08CRCNODsHN0FVMRF#sRHDMoCFR#kCsOR#8CHIoMN
sCNs00H0LkC$R#Mk_LHHD0Mk_8R#:R0MsHoN;
0H0sLCk0RM#$_HLkDM0H_R8kF7VRWb_V_8N8#RkL:MRC0$H0RRH#"NIC	
";
M
C8WR7__VbN#88k
L;
ONsECH0Os0kC0RsDVRFR_7WVNb_8k8#L#RH
-
-R0N0skHL08CRCNODsHN0FVMRF#sRHDMoCFR#kCsOR#8CHIoMNRsC
0N0skHL0#CR$LM_k0HDH8M_kRR:#H0sM
o;Ns00H0LkC$R#Mk_LHHD0Mk_8RRFVsR0D:sRNO0EHCkO0sHCR#IR"C"N	;-

-FRwsHR#MCoDRk#FsROC7RW,NEsOHO0C0CksRF#EkRD8L8CRk$ll
0N0skHL0#CR$LM_D	NO_GLFRL:RFCFDN
M;Ns00H0LkC$R#MD_LN_O	LRFGFsVR0:DRRONsECH0Os0kC#RHRk0sC
;
LHCoMC

Ms8R0
D;
-
--------------------------------------------------------------------------------------
-
DsHLNRs$Q   ,q7W)
 ;kR#CQ   38#0_oDFH4O_43ncN;DD
Ck#Rq7W)7 3WF_wkNM80MHF_lOFbD3ND
;
CHM007$RWb_V_P8HR
H#
MoCCOsHR#5
HIo_HE80Ru:Rma1QQRe :.=RdC;
GIb_HE80Ru:Rma1QQRe :U=R;C
HCOC_FDlbHONMCRR:Q hatR ):j=R;N
VHV0EksD_F8kMRQ:Rhta  :)R=
Rj2
;
b0FsRN5
RH:RM0R#8F_Do_HOP0COF#s5HIo_HE80RC+RGIb_HE80RI8FMR0Fj
2;LRR:H#MR0D8_FOoH_OPC05Fs#_HoI0H8ERR+C_GbI0H8EFR8IFM0R;j2
8sMRH:RM0R#8F_Do_HOP0COF.s5RI8FMR0Fj
2;xF:Rk#0R0D8_FOoH_OPC05Fs#_HoI0H8ERR+C_GbI0H8EFR8IFM0R;j2
N#00:k#R0FkR8#0_oDFHPO_CFO0sR5(8MFI0jFR2;
2
-
-R0N0skHL08CRCNODsHN0FVMRF#sRHDMoCFR#kCsOR#8CHIoMN
sCNs00H0LkC$R#Mk_LHHD0Mk_8R#:R0MsHoN;
0H0sLCk0RM#$_HLkDM0H_R8kF7VRWb_V_P8HRC:RM00H$#RHRC"IN;	"
M
C8WR7__Vb8;HP
N

sHOE00COkRsCsR0DF7VRWb_V_P8HR
H#
R--Ns00H0LkCCR8OsDNNF0HMFRVsHR#MCoDRk#FsROC8HC#oNMIs
CRNs00H0LkC$R#Mk_LHHD0Mk_8R#:R0MsHoN;
0H0sLCk0RM#$_HLkDM0H_R8kFsVR0:DRRONsECH0Os0kC#RHRC"IN;	"
-
-RswFRM#HoRDC#sFkO7CRWN,RsHOE00COkRsC#kEFDL8RCkR8l
l$Ns00H0LkC$R#MD_LN_O	LRFG:FRLFNDCMN;
0H0sLCk0RM#$_NLDOL	_FFGRV0RsDRR:NEsOHO0C0CksRRH#0Csk;L

CMoH
C

Ms8R0
D;
--------------------------------------------------------------------------------------------
-
DsHLNRs$Q   ,q7W)
 ;kR#CQ   38#0_oDFH4O_43ncN;DD
Ck#Rq7W)7 3WF_wkNM80MHF_lOFbD3ND
;
CHM007$RWb_V_0VD.HHR#o

CsMCH5OR
o#H_8IH0:ERR1umQeaQ =R:R;.d
bCG_8IH0:ERR1umQeaQ =R:R
U;Hx#HCRR:Q hatR ):d=R.;
2
F
bs50R
:NRRRHM#_08DHFoOC_POs0F5o#H_8IH0+ERRGRCbH_I8R0E8MFI0jFR2s;
M:8RRRHM#_08DHFoOC_POs0F58.RF0IMF2Rj;:
xR0FkR8#0_oDFHPO_CFO0s#5HH-xC4FR8IFM0R;j2
N#00:k#R0FkR8#0_oDFHPO_CFO0sR5(8MFI0jFR2;
2
-
-R0N0skHL08CRCNODsHN0FVMRF#sRHDMoCFR#kCsOR#8CHIoMN
sCNs00H0LkC$R#Mk_LHHD0Mk_8R#:R0MsHoN;
0H0sLCk0RM#$_HLkDM0H_R8kF7VRWb_V_0VD.:HRR0CMHR0$H"#RI	CN"
;

8CMR_7WVVb_DH0.;N

sHOE00COkRsCsR0DF7VRWb_V_0VD.HHR#-

-0RN0LsHkR0C8DCON0sNHRFMVRFs#oHMD#CRFOksCCR8#MHoICNsR0
N0LsHkR0C#_$MLDkH0_HM8:kRRs#0H;Mo
0N0skHL0#CR$LM_k0HDH8M_kVRFRDs0RN:RsHOE00COkRsCH"#RI	CN"
;
-w-RF#sRHDMoCFR#kCsOR,7WRONsECH0Os0kCER#F8kDRRLC8lkl$0
N0LsHkR0C#_$MLODN	F_LGRR:LDFFC;NM
0N0skHL0#CR$LM_D	NO_GLFRRFVsR0D:sRNO0EHCkO0sHCR#sR0k
C;
oLCH
M
CRM8s;0D
-

-----------------------------------------------------------------------------------------
--
LDHs$NsR Q  W,7q;) 
Ck#R Q  03#8F_Do_HO4c4n3DND;#
kCWR7q3) 7wW_F8kMNF0HMF_OlNb3D
D;
0CMHR0$7VW_b._HVRD0H
#
oCCMsRHO5H
#oH_I8R0E:mRu1QQae: R=dR.;G
CbH_I8R0E:mRu1QQae: R=;RU
HH#x:CRR1umQeaQ =R:R;d.
HH#o:MRRaQh )t RR:=4;
2
F
bs50R
:NRRRHM#_08DHFoOC_POs0F5HH#x4C-RI8FMR0Fj
2;sRM8:MRHR8#0_oDFHPO_CFO0sR5.8MFI0jFR2x;
:kRF00R#8F_Do_HOP0COF#s5HIo_HE80RC+RGIb_HE80RI8FMR0Fj
2;#00NkR#:FRk0#_08DHFoOC_POs0F58(RF0IMF2Rj

2;
R--Ns00H0LkCCR8OsDNNF0HMFRVsHR#MCoDRk#FsROC8HC#oNMIsNC
0H0sLCk0RM#$_HLkDM0H_R8k:0R#soHM;0
N0LsHkR0C#_$MLDkH0_HM8FkRVWR7__VbHD.V0RR:CHM00H$R#IR"C"N	;C

M78RWb_V_VH.D
0;
ONsECH0Os0kC0RsDVRFR_7WVHb_.0VDR
H#
R--Ns00H0LkCCR8OsDNNF0HMFRVsHR#MCoDRk#FsROC8HC#oNMIs
CRNs00H0LkC$R#Mk_LHHD0Mk_8R#:R0MsHoN;
0H0sLCk0RM#$_HLkDM0H_R8kFsVR0:DRRONsECH0Os0kC#RHRC"IN;	"
-
-RswFRM#HoRDC#sFkO7CRWN,RsHOE00COkRsC#kEFDL8RCkR8l
l$Ns00H0LkC$R#MD_LN_O	LRFG:FRLFNDCMN;
0H0sLCk0RM#$_NLDOL	_FFGRV0RsDRR:NEsOHO0C0CksRRH#0Csk;L

CMoH
M
C80RsD
;
---------------------------------------------------------------------------------------------
--
LDHs$NsR Q  W,7q;) 
Ck#R Q  03#8F_Do_HO4c4n3DND;#
kCWR7q3) 7wW_F8kMNF0HMF_OlNb3D
D;
0CMHR0$7VW_bk_lDH0R#o

CsMCH5OR
o#H_8IH0:ERR1umQeaQ =R:R;.d
bCG_8IH0:ERR1umQeaQ =R:R
U;HCCC_lOFbNDHMROC:hRQa  t)=R:R2j
;b

FRs05R
N:MRHR8#0_oDFHPO_CFO0sH5#oH_I8R0E+GRCbH_I8R0E8MFI0jFR2L;
RH:RM0R#8F_Do_HOP0COF#s5HIo_HE80RC+RGIb_HE80RI8FMR0Fj
2;sRM8:MRHR8#0_oDFHPO_CFO0sR5.8MFI0jFR2x;
:kRF00R#8F_Do_HOP0COF#s5HIo_HE80RC+RGIb_HE80RI8FMR0Fj
2;#00NkR#:FRk0#_08DHFoOC_POs0F58(RF0IMF2Rj

2;
R--Ns00H0LkCCR8OsDNNF0HMFRVsHR#MCoDRk#FsROC8HC#oNMIsNC
0H0sLCk0RM#$_HLkDM0H_R8k:0R#soHM;0
N0LsHkR0C#_$MLDkH0_HM8FkRVWR7__Vbl0kDRC:RM00H$#RHRC"IN;	"
M
C8WR7__Vbl0kD;N

sHOE00COkRsCsR0DF7VRWb_V_Dlk0#RH
-
-R0N0skHL08CRCNODsHN0FVMRF#sRHDMoCFR#kCsOR#8CHIoMNRsC
0N0skHL0#CR$LM_k0HDH8M_kRR:#H0sM
o;Ns00H0LkC$R#Mk_LHHD0Mk_8RRFVsR0D:sRNO0EHCkO0sHCR#IR"C"N	;-

-FRwsHR#MCoDRk#FsROC7RW,NEsOHO0C0CksRF#EkRD8L8CRk$ll
0N0skHL0#CR$LM_D	NO_GLFRL:RFCFDN
M;Ns00H0LkC$R#MD_LN_O	LRFGFsVR0:DRRONsECH0Os0kC#RHRk0sC
;
LHCoM


CRM8s;0D
-

---------------------------------------------------------------------------------------------D

HNLssQ$R ,  Rq7W)
 ;kR#CQ   38#0_oDFH4O_43ncN;DD
Ck#Rq7W)7 3WF_wkNM80MHF_lOFbs_NH30EN;DD
M
C0$H0R_7WH_MOo$sNR
H#
MoCCOsHRH5I8R0E:FRb#HH0P:CR=2RU;b

FRs05:NRRRHM#_08DHFoOC_POs0F58IH04E-RI8FMR0Fj
2;O:HRRRHM#_08DHFoOx;
:kRF00R#8F_Do_HOP0COFIs5HE80-84RF0IMF2Rj2
;
-N-R0H0sLCk0RO8CDNNs0MHFRsVFRM#HoRDC#sFkO8CRCo#HMsINC0
N0LsHkR0C#_$MLDkH0_HM8:kRRs#0H;Mo
0N0skHL0#CR$LM_k0HDH8M_kVRFR_7WH_MOo$sNRC:RM00H$#RHRC"IN;	"
M
C8WR7_OHM_Nos$
;

ONsECH0Os0kC0RsDVRFR_7WH_MOo$sNR
H#
R--Ns00H0LkCCR8OsDNNF0HMFRVsHR#MCoDRk#FsROC8HC#oNMIs
CRNs00H0LkC$R#Mk_LHHD0Mk_8R#:R0MsHoN;
0H0sLCk0RM#$_HLkDM0H_R8kFsVR0:DRRONsECH0Os0kC#RHRC"IN;	"
-
-RswFRM#HoRDC#sFkO7CRWN,RsHOE00COkRsC#kEFDL8RCkR8l
l$Ns00H0LkC$R#MD_LN_O	LRFG:FRLFNDCMN;
0H0sLCk0RM#$_NLDOL	_FFGRV0RsDRR:NEsOHO0C0CksRRH#0Csk;


LHCoMC

Ms8R0
D;
-
------------------------------------------------------------------------------------------
--
LDHs$NsR Q  W,7q;) 
Ck#R Q  03#8F_Do_HO4c4n3DND;#
kCWR7q3) 7NWbOo	NCN#3D
D;kR#C7)Wq I38_kVFM08NH_FMObFl3DND;C

M00H$WR7_#DLE#RH
C
oMHCsO
R5qH_I8R0E:mRu1QQae: R=;RU
_1]I0H8ERR:uQm1a QeRR:=d;
2
F
bs50R
:qRRRHM#_08DHFoOC_POs0F5Iq_HE80-84RF0IMF2Rj;]
1RH:RM0R#8F_Do_HOP0COF1s5]H_I8-0E4FR8IFM0R;j2
_1]a:BRRRHM#_08DHFoOA;
:kRF00R#8F_Do_HOP0COFqs5_8IH04E-RI8FMR0Fj22
;-

-0RN0LsHkR0C8DCON0sNHRFMVRFs#oHMD#CRFOksCCR8#MHoICNs
0N0skHL0#CR$LM_k0HDH8M_kRR:#H0sM
o;Ns00H0LkC$R#Mk_LHHD0Mk_8RRFV7DW_LR#E:MRC0$H0RRH#"NIC	
";
M
C8WR7_#DLE
;
NEsOHO0C0CksRDs0RRFV7DW_LR#EH
#
-N-R0H0sLCk0RO8CDNNs0MHFRsVFRM#HoRDC#sFkO8CRCo#HMsINCNR
0H0sLCk0RM#$_HLkDM0H_R8k:0R#soHM;0
N0LsHkR0C#_$MLDkH0_HM8FkRV0RsDRR:NEsOHO0C0CksRRH#"NIC	
";
R--wRFs#oHMD#CRFOksCWR7,sRNO0EHCkO0s#CREDFk8CRLRl8klN$
0H0sLCk0RM#$_NLDOL	_F:GRRFLFDMCN;0
N0LsHkR0C#_$MLODN	F_LGVRFRDs0RN:RsHOE00COkRsCH0#Rs;kC
L

CMoH
M
C80RsD
;

--------------------------------------------------------------------------------------------
-
DsHLNRs$Q   ,q7W)
 ;kR#CQ   38#0_oDFH4O_43ncN;DD
Ck#Rq7W)7 3WF_wkNM80MHF_lOFbD3NDk;
#7CRW q)3b7WNNO	o3C#N;DD
M
C0$H0R_7WDRx8H
#
oCCMsRHO5_
NI0H8ERR:uQm1a QeRR:=U;
2
F
bs50R
:NRRRHM#_08DHFoOC_POs0F5IN_HE80-84RF0IMF2Rj;C
8ORR:FRk0#_08DHFoOC_POs0F5IN_HE80-84RF0IMF2Rj;M
CORR:FRk0#_08DHFoOC_POs0F50LH_8IH0NE5_8IH0RE28MFI0jFR2;
2
-
-R0N0skHL08CRCNODsHN0FVMRF#sRHDMoCFR#kCsOR#8CHIoMN
sCNs00H0LkC$R#Mk_LHHD0Mk_8R#:R0MsHoN;
0H0sLCk0RM#$_HLkDM0H_R8kF7VRWx_D8RR:CHM00H$R#IR"C"N	;C

M78RWx_D8
;

ONsECH0Os0kC0RsDVRFR_7WDRx8H
#
-N-R0H0sLCk0RO8CDNNs0MHFRsVFRM#HoRDC#sFkO8CRCo#HMsINCNR
0H0sLCk0RM#$_HLkDM0H_R8k:0R#soHM;0
N0LsHkR0C#_$MLDkH0_HM8FkRV0RsDRR:NEsOHO0C0CksRRH#"NIC	
";
R--wRFs#oHMD#CRFOksCWR7,sRNO0EHCkO0s#CREDFk8CRLRl8klN$
0H0sLCk0RM#$_NLDOL	_F:GRRFLFDMCN;0
N0LsHkR0C#_$MLODN	F_LGVRFRDs0RN:RsHOE00COkRsCH0#Rs;kC
L

CMoH
M
C80RsD
;

-------------------------------------------------------------------------------------------
H
DLssN$ RQ 7 ,W q);#
kC RQ # 30D8_FOoH_n44cD3NDk;
#7CRW q)3b7WNNO	o3C#N;DD
Ck#Rq7W)8 3IF_VkNM80MHF_lOFbD3ND
;
CHM007$RWN_s#HER#o

CsMCH5OR
Iq_HE80Ru:Rma1QQRe :U=R;]
1_8IH0:ERR1umQeaQ =R:R2d
;b

FRs05R
q:MRHR8#0_oDFHPO_CFO0s_5qI0H8ER-48MFI0jFR27;
q_aqa:BRRRHM#_08DHFoO1;
]RR:H#MR0D8_FOoH_OPC05Fs1I]_HE80-84RF0IMF2Rj;]
1_RaB:MRHR8#0_oDFH
O;ARR:FRk0#_08DHFoOC_POs0F5Iq_HE80-84RF0IMF2Rj

2;
R--Ns00H0LkCCR8OsDNNF0HMFRVsHR#MCoDRk#FsROC8HC#oNMIsNC
0H0sLCk0RM#$_HLkDM0H_R8k:0R#soHM;0
N0LsHkR0C#_$MLDkH0_HM8FkRVWR7_#sNERR:CHM00H$R#IR"C"N	;


CRM87sW_N;#E
s
NO0EHCkO0ssCR0FDRVWR7_#sNE#RH
-
-R0N0skHL08CRCNODsHN0FVMRF#sRHDMoCFR#kCsOR#8CHIoMNRsC
0N0skHL0#CR$LM_k0HDH8M_kRR:#H0sM
o;Ns00H0LkC$R#Mk_LHHD0Mk_8RRFVsR0D:sRNO0EHCkO0sHCR#IR"C"N	;-

-FRwsHR#MCoDRk#FsROC7RW,NEsOHO0C0CksRF#EkRD8L8CRk$ll
0N0skHL0#CR$LM_D	NO_GLFRL:RFCFDN
M;Ns00H0LkC$R#MD_LN_O	LRFGFsVR0:DRRONsECH0Os0kC#RHRk0sC
;
LHCoMC

Ms8R0
D;
-
--------------------------------------------------------------------------------------
-
DsHLNRs$Q   ,q7W)
 ;kR#CQ   38#0_oDFH4O_43ncN;DD
Ck#Rq7W)7 3WObN	CNo#D3NDk;
#7CRW q)3_8IVMFk8HN0FOM_F3lbN;DD
M
C0$H0R_7WsEL#R
H#
MoCCOsHRq5
_8IH0:ERR1umQeaQ =R:R
U;1I]_HE80Ru:Rma1QQRe :d=R

2;
sbF0
R5qRR:H#MR0D8_FOoH_OPC05FsqH_I8-0E4FR8IFM0R;j2
R1]:MRHR8#0_oDFHPO_CFO0s]51_8IH04E-RI8FMR0Fj
2;1a]_BRR:H#MR0D8_FOoH;:
AR0FkR8#0_oDFHPO_CFO0s_5qI0H8ER-48MFI0jFR2;
2
-
-R0N0skHL08CRCNODsHN0FVMRF#sRHDMoCFR#kCsOR#8CHIoMN
sCNs00H0LkC$R#Mk_LHHD0Mk_8R#:R0MsHoN;
0H0sLCk0RM#$_HLkDM0H_R8kF7VRWL_s#:ERR0CMHR0$H"#RI	CN"
;
CRM87sW_L;#E
s
NO0EHCkO0ssCR0FDRVWR7_#sLE#RH
-
-R0N0skHL08CRCNODsHN0FVMRF#sRHDMoCFR#kCsOR#8CHIoMNRsC
0N0skHL0#CR$LM_k0HDH8M_kRR:#H0sM
o;Ns00H0LkC$R#Mk_LHHD0Mk_8RRFVsR0D:sRNO0EHCkO0sHCR#IR"C"N	;-

-FRwsHR#MCoDRk#FsROC7RW,NEsOHO0C0CksRF#EkRD8L8CRk$ll
0N0skHL0#CR$LM_D	NO_GLFRL:RFCFDN
M;Ns00H0LkC$R#MD_LN_O	LRFGFsVR0:DRRONsECH0Os0kC#RHRk0sC
;
LHCoMC

Ms8R0
D;
-

------------------------------------------------------------------------------------------------
LDHs$NsR Q  W,7q;) 
Ck#R Q  03#8F_Do_HO4c4n3DND;#
kCWR7q3) 7wW_F8kMNF0HMF_OlNb_sEH03DND;C

M00H$WR7_0OMss_oNH$R#C
oMHCsOIR5HE80Ru:Rma1QQRe :U=R2
;
b0FsRD5O	RR:H#MR0D8_FOoH;R
RRRRRs_#0MRR:H#MR0D8_FOoH;R
RRRRRH0MH_:MRRRHM#_08DHFoOR;
RRRRRNDF8R_M:MRHR8#0_oDFH
O;RRRRRNR80:NRRRHM#_08DHFoOC_POs0F58IH04E-RI8FMR0Fj
2;RRRRRCROMRR:H#MR0D8_FOoH;R
RRRRROMFk0RR:FRk0#_08DHFoOC_POs0F58IH04E-RI8FMR0Fj;22



-N-R0H0sLCk0RO8CDNNs0MHFRsVFRM#HoRDC#sFkO8CRCo#HMsINC0
N0LsHkR0C#_$MLDkH0_HM8:kRRs#0H;Mo
0N0skHL0#CR$LM_k0HDH8M_kVRFR_7WOsM0_Nos$RR:CHM00H$R#IR"C"N	;C

M78RWM_O0os_s;N$
N

sHOE00COkRsCsR0DF7VRWM_O0os_sRN$H
#
-N-R0H0sLCk0RO8CDNNs0MHFRsVFRM#HoRDC#sFkO8CRCo#HMsINCNR
0H0sLCk0RM#$_HLkDM0H_R8k:0R#soHM;0
N0LsHkR0C#_$MLDkH0_HM8FkRV0RsDRR:NEsOHO0C0CksRRH#"NIC	
";
R--wRFs#oHMD#CRFOksCWR7,sRNO0EHCkO0s#CREDFk8CRLRl8klN$
0H0sLCk0RM#$_NLDOL	_F:GRRFLFDMCN;0
N0LsHkR0C#_$MLODN	F_LGVRFRDs0RN:RsHOE00COkRsCH0#Rs;kC
C
Lo
HM
8CMRDs0;



-
--------------------------------------------------------------------------------------------------H
DLssN$ RQ 7 ,W q);#
kC RQ # 30D8_FOoH_n44cD3NDk;
#7CRW q)3_7WwMFk8HN0FOM_F_lbN0sHED3ND
;
CHM007$RWs_oNL$.HHMR#C
oMHCsOIR5HE80Ru:Rma1QQRe :U=R2
;
b0FsRR5o:MRHR8#0_oDFHPO_CFO0sH5I8-0E4FR8IFM0R;j2
RRRRLRRRF:Rk#0R0D8_FOoH_OPC05FsI0H8ER-48MFI0jFR2
2;
R--Ns00H0LkCCR8OsDNNF0HMFRVsHR#MCoDRk#FsROC8HC#oNMIsRC
RRRRRNRR0H0sLCk0RM#$_HLkDM0H_R8k:0R#soHM;R
RRRRRR0RN0LsHkR0C#_$MLDkH0_HM8FkRVWR7_Nos$H.LMRR:CHM00H$R#IR"C"N	;C

M78RWs_oNL$.H
M;
s
NO0EHCkO0ssCR0FDRVWR7_Nos$H.LM#RH
-
-R0N0skHL08CRCNODsHN0FVMRF#sRHDMoCFR#kCsOR#8CHIoMNRsC
0N0skHL0#CR$LM_k0HDH8M_kRR:#H0sM
o;Ns00H0LkC$R#Mk_LHHD0Mk_8RRFVsR0D:sRNO0EHCkO0sHCR#IR"C"N	;-

-FRwsHR#MCoDRk#FsROC7RW,NEsOHO0C0CksRF#EkRD8L8CRk$ll
0N0skHL0#CR$LM_D	NO_GLFRL:RFCFDN
M;Ns00H0LkC$R#MD_LN_O	LRFGFsVR0:DRRONsECH0Os0kC#RHRk0sC
;
LHCoMC

Ms8R0
D;
---------------------------------------------------------------------------------------------------
D

HNLssQ$R ,  7)Wq k;
#QCR 3  #_08DHFoO4_4nNc3D
D;kR#C7)Wq W37_kwFM08NH_FMObFl_HNs0NE3D
D;
0CMHR0$7LW_HoM.sRN$Ho#
CsMCH5ORI0H8ERR:uQm1a QeRR:=U
2;
sbF0LR5RH:RM0R#8F_Do_HOP0COFIs5HE80-84RF0IMF2Rj;R
RRRRRoRR:FRk0#_08DHFoOC_POs0F58IH04E-RI8FMR0Fj;22
-
-R0N0skHL08CRCNODsHN0FVMRF#sRHDMoCFR#kCsOR#8CHIoMN
sCRRRRRRRRNs00H0LkC$R#Mk_LHHD0Mk_8R#:R0MsHoR;
RRRRRNRR0H0sLCk0RM#$_HLkDM0H_R8kF7VRWH_LMs.oN:$RR0CMHR0$H"#RI	CN"
;
CRM87LW_HoM.s;N$
N

sHOE00COkRsCsR0DF7VRWH_LMs.oNH$R#-

-0RN0LsHkR0C8DCON0sNHRFMVRFs#oHMD#CRFOksCCR8#MHoICNsR0
N0LsHkR0C#_$MLDkH0_HM8:kRRs#0H;Mo
0N0skHL0#CR$LM_k0HDH8M_kVRFRDs0RN:RsHOE00COkRsCH"#RI	CN"
;
-w-RF#sRHDMoCFR#kCsOR,7WRONsECH0Os0kCER#F8kDRRLC8lkl$0
N0LsHkR0C#_$MLODN	F_LGRR:LDFFC;NM
0N0skHL0#CR$LM_D	NO_GLFRRFVsR0D:sRNO0EHCkO0sHCR#sR0k
C;
oLCH
M
CRM8s;0D
-

-------------------------------------------------------------------------------------------------
-

H
DLssN$ RQ R ,7)Wq k;
#QCR 3  #_08DHFoO4_4nNc3D
D;kR#C7)Wq W37_kwFM08NH_FMObFl_HNs0NE3D
D;
0CMHR0$78W_HbP_HRbCHo#
CsMCH5ORNH_I8R0E:mRu1QQae: R=;RURIL_HE80Ru:Rma1QQRe :U=R;O
0_8lFCRR:hzqa)Rqp:j=R;CRslF_l8:CRRahqzp)qRR:=4M;
k#l_0CNo#RR:uQm1a QeRR:=.#;R0DND_8lFCRR:hzqa)Rqp:4=R;#
s0F_l8:CRRahqzp)qRR:=4;R2
F
bs50RORD	:MRHR8#0_oDFH
O;s_#0MRR:H#MR0D8_FOoH;M
CRH:RM0R#8F_Do;HO
:NRRRHM#_08DHFoOC_POs0F5IN_HE80-84RF0IMF2Rj;R
L:MRHR8#0_oDFHPO_CFO0s_5LI0H8ER-48MFI0jFR2J;
kHF0CRM0:kRF00R#8F_Do_HOP0COFNs5_8IH04E-RI8FMR0Fj
2;sNClHCM8sRR:FRk0#_08DHFoOC_POs0F5IL_HE80-84RF0IMF2Rj;H
8PCH8__L$jRR:FRk0#_08DHFoO;R2
-
-R0N0skHL08CRCNODsHN0FVMRF#sRHDMoCFR#kCsOR#8CHIoMN
sCRRRRRRRRNs00H0LkC$R#Mk_LHHD0Mk_8R#:R0MsHoR;
RRRRRNRR0H0sLCk0RM#$_HLkDM0H_R8kF7VRWH_8PH_bb:CRR0CMHR0$H"#RI	CN"
;

8CMR_7W8_HPbCHb;


NEsOHO0C0CksRDs0RRFV78W_HbP_HRbCH
#
-N-R0H0sLCk0RO8CDNNs0MHFRsVFRM#HoRDC#sFkO8CRCo#HMsINCNR
0H0sLCk0RM#$_HLkDM0H_R8k:0R#soHM;0
N0LsHkR0C#_$MLDkH0_HM8FkRV0RsDRR:NEsOHO0C0CksRRH#"NIC	
";
R--wRFs#oHMD#CRFOksCWR7,sRNO0EHCkO0s#CREDFk8CRLRl8klN$
0H0sLCk0RM#$_NLDOL	_F:GRRFLFDMCN;0
N0LsHkR0C#_$MLODN	F_LGVRFRDs0RN:RsHOE00COkRsCH0#Rs;kC
C
Lo
HM
M
C80RsD
;

------------------------------------------------------------------------------------------------
--DsHLNRs$Q   ,q7W)
 ;kR#CQ   38#0_oDFH4O_43ncN;DD
Ck#Rq7W)7 3WF_wkNM80MHF_lOFbs_NH30EN;DD
M
C0$H0R_7W#0Js_bbHC#RH
MoCCOsHRH5I8R0E:mRu1QQae: R=;R.R_0OlCF8Rh:Rq)azq:pR=;Rj
lMk_N#0oRC#:mRu1QQae: R=;R.RN#0DlD_FR8C:qRhaqz)p=R:R
4;s_#0lCF8Rh:Rq)azq:pR=RR42
;
b0FsRD5O	RR:H#MR0D8_FOoH;#
s0R_M:MRHR8#0_oDFH
O;C:MRRRHM#_08DHFoON;
RH:RM0R#8F_Do_HOP0COFIs5HE80-84RF0IMF2Rj;F
sF:0RR0FkR8#0_oDFHPO_CFO0sI55HE80+/42.R-48MFI0jFR2;R2
-
-R0N0skHL08CRCNODsHN0FVMRF#sRHDMoCFR#kCsOR#8CHIoMN
sCRRRRRRRRNs00H0LkC$R#Mk_LHHD0Mk_8R#:R0MsHoR;
RRRRRNRR0H0sLCk0RM#$_HLkDM0H_R8kF7VRWJ_#sb0_HRbC:MRC0$H0RRH#"NIC	
";
8CMR_7W#0Js_bbHC
;

ONsECH0Os0kC0RsDVRFR_7W#0Js_bbHC#RH
-
-R0N0skHL08CRCNODsHN0FVMRF#sRHDMoCFR#kCsOR#8CHIoMNRsC
0N0skHL0#CR$LM_k0HDH8M_kRR:#H0sM
o;Ns00H0LkC$R#Mk_LHHD0Mk_8RRFVsR0D:sRNO0EHCkO0sHCR#IR"C"N	;-

-FRwsHR#MCoDRk#FsROC7RW,NEsOHO0C0CksRF#EkRD8L8CRk$ll
0N0skHL0#CR$LM_D	NO_GLFRL:RFCFDN
M;Ns00H0LkC$R#MD_LN_O	LRFGFsVR0:DRRONsECH0Os0kC#RHRk0sC
;
LHCoMC

Ms8R0
D;
-
--------------------------------------------------------------------------------------------------D

HNLssQ$R ,  7)Wq k;
#QCR 3  #_08DHFoO4_4nNc3D
D;kR#C7)Wq W37_kwFM08NH_FMObFl_HNs0NE3D
D;
0CMHR0$7lW_k_D0bCHbR
H#oCCMsRHO5_
NI0H8ERR:uQm1a QeRR:=U
;RLH_I8R0E:mRu1QQae: R=;RU
lMk_N#0oRC#:mRu1QQae: R=;R.R0
#N_DDlCF8Rh:Rq)azq:pR=;R4
0s#_8lFCRR:hzqa)Rqp:4=R
RRRRRRRR
2;
sbF0
R5ORD	:MRHR8#0_oDFHRO;
0s#_:MRRRHM#_08DHFoOC;
MRR:H#MR0D8_FOoH;0R
ORR:H#MR0D8_FOoH;R
N:MRHR8#0_oDFHPO_CFO0s_5NI0H8ER-48MFI0jFR2L;
RH:RM0R#8F_Do_HOP0COFLs5_8IH04E-RI8FMR0Fj
2;b8sFkRO0:kRF00R#8F_Do_HOP0COFNs5_8IH0+ERRIL_HE80-84RF0IMF2Rj

2;
R--Ns00H0LkCCR8OsDNNF0HMFRVsHR#MCoDRk#FsROC8HC#oNMIsRC
RRRRRNRR0H0sLCk0RM#$_HLkDM0H_R8k:0R#soHM;R
RRRRRR0RN0LsHkR0C#_$MLDkH0_HM8FkRVWR7_Dlk0H_bb:CRR0CMHR0$H"#RI	CN"
;
CRM87lW_k_D0bCHb;N

sHOE00COkRsCsR0DF7VRWk_lDb0_HRbCH
#
-N-R0H0sLCk0RO8CDNNs0MHFRsVFRM#HoRDC#sFkO8CRCo#HMsINCNR
0H0sLCk0RM#$_HLkDM0H_R8k:0R#soHM;0
N0LsHkR0C#_$MLDkH0_HM8FkRV0RsDRR:NEsOHO0C0CksRRH#"NIC	
";
R--wRFs#oHMD#CRFOksCWR7,sRNO0EHCkO0s#CREDFk8CRLRl8klN$
0H0sLCk0RM#$_NLDOL	_F:GRRFLFDMCN;0
N0LsHkR0C#_$MLODN	F_LGVRFRDs0RN:RsHOE00COkRsCH0#Rs;kC
C
Lo
HM
M
C80RsD
;
------------------------------------------------------------------------------------
H
DLssN$ RQ 7 ,W q);#
kC RQ # 30D8_FOoH_n44cD3NDk;
#7CRW q)3b7WNNO	o3C#N;DD
Ck#Rq7W)7 3WF_wkNM80MHF_lOFbs_NH30EN;DD
M
C0$H0R_7Wb8sF_l#k_bbHC#RH
C
oMHCsO
R5NH_I8R0E:mRu1QQae: R=;R.
IL_HE80Ru:Rma1QQRe :.=R;k
MlM_Hb#k0Ru:Rma1QQRe :.=R;k
#lH_I8R0E:mRu1QQae: R=;Rc
lMk_N#0oRC#:mRu1QQae: R=;R.
N#0DlD_FR8C:qRhaqz)p=R:R
4;s_#0lCF8Rh:Rq)azq:pR=RR4

2;
sbF0
R5
	ODRH:RM0R#8F_Do;HO
0s#_:MRRRHM#_08DHFoOC;
MRR:H#MR0D8_FOoH;O
0RH:RM0R#8F_Do;HO
:NRRRHM#_08DHFoOC_POs0F5IN_HE80*lMk_bHMk-0#4FR8IFM0R;j2
:LRRRHM#_08DHFoOC_POs0F5IL_HE80*lMk_bHMk-0#4FR8IFM0R;j2
l#kRF:Rk#0R0D8_FOoH_OPC05Fs#_klI0H8ER-48MFI0jFR2;R2
-
-R0N0skHL08CRCNODsHN0FVMRF#sRHDMoCFR#kCsOR#8CHIoMN
sCRRRRRRRRNs00H0LkC$R#Mk_LHHD0Mk_8R#:R0MsHoR;
RRRRRNRR0H0sLCk0RM#$_HLkDM0H_R8kF7VRWs_bF#8_kbl_HRbC:MRC0$H0RRH#"NIC	
";
8CMR_7Wb8sF_l#k_bbHC
;
NEsOHO0C0CksRDs0RRFV7bW_s_F8#_klbCHbR
H#
R--Ns00H0LkCCR8OsDNNF0HMFRVsHR#MCoDRk#FsROC8HC#oNMIs
CRNs00H0LkC$R#Mk_LHHD0Mk_8R#:R0MsHoN;
0H0sLCk0RM#$_HLkDM0H_R8kFsVR0:DRRONsECH0Os0kC#RHRC"IN;	"
-
-RswFRM#HoRDC#sFkO7CRWN,RsHOE00COkRsC#kEFDL8RCkR8l
l$Ns00H0LkC$R#MD_LN_O	LRFG:FRLFNDCMN;
0H0sLCk0RM#$_NLDOL	_FFGRV0RsDRR:NEsOHO0C0CksRRH#0Csk;L

CMoH
M
C80RsD
;

----------------------------------------------------------------------------D

HNLssQ$R ,  7)Wq k;
#QCR 3  #_08DHFoO4_4nNc3D
D;kR#C7)Wq W37_kwFM08NH_FMObFl_HNs0NE3D
D;
0CMHR0$7LW_OR_UHb#
FRs05bON0Cks_	ODRH:RM0R#8F_Do;HO
8kbN_0CORD	:MRHR8#0_oDFH
O;O0Nbk_sCC:MRRRHM#_08DHFoOk;
b08NCM_CRH:RM0R#8F_Do;HO
H#EV80_sRR:H#MR0D8_FOoH;F
l8:CRRRHM#_08DHFoO#;
HRR:H#MR0D8_FOoH;H
bMM_HbRk0:MRHR8#0_oDFH
O;Fbk0k80_NR0N:MRHR8#0_oDFH
O;HHO_M0bkRF:Rk#0R0D8_FOoH;N
80FN_k:0RR0FkR8#0_oDFH
O;#:FRR0FkR8#0_oDFH2OR;-

-0RN0LsHkR0C8DCON0sNHRFMVRFs#oHMD#CRFOksCCR8#MHoICNs
RRRRRRRR0N0skHL0#CR$LM_k0HDH8M_kRR:#H0sM
o;RRRRRRRRNs00H0LkC$R#Mk_LHHD0Mk_8RRFV7LW_OR_U:MRC0$H0RRH#"NIC	
";
M
C8WR7__LOU
;
NEsOHO0C0CksRDs0RRFV7LW_OR_UH
#
-N-R0H0sLCk0RO8CDNNs0MHFRsVFRM#HoRDC#sFkO8CRCo#HMsINCNR
0H0sLCk0RM#$_HLkDM0H_R8k:0R#soHM;0
N0LsHkR0C#_$MLDkH0_HM8FkRV0RsDRR:NEsOHO0C0CksRRH#"NIC	
";R-
-RswFRM#HoRDC#sFkO7CRWN,RsHOE00COkRsC#kEFDL8RCkR8l
l$Ns00H0LkC$R#MD_LN_O	LRFG:FRLFNDCMN;
0H0sLCk0RM#$_NLDOL	_FFGRV0RsDRR:NEsOHO0C0CksRRH#0Csk;


LHCoMM
C80RsD
;
---------------------------------------------------------------------------------
--
H
DLssN$ RQ 7 ,W q);#
kC RQ # 30D8_FOoH_n44cD3NDk;
#7CRW q)3_7WwMFk8HN0FOM_F_lbN0sHED3ND
;
CHM007$RWO_L_HgR#F
bs50RO0Nbk_sCORD	:MRHR8#0_oDFH
O;kNb80OC_D:	RRRHM#_08DHFoOO;
Nkb0sCC_MRR:H#MR0D8_FOoH;b
k8CN0_RCM:MRHR8#0_oDFH
O;#VEH0s_8RH:RM0R#8F_Do;HO
8lFC:4RRRHM#_08DHFoOl;
F.8CRH:RM0R#8F_Do;HO
R#H:MRHR8#0_oDFH
O;b_HMHkMb0RR:H#MR0D8_FOoH;k
F00bk_08NNRR:H#MR0D8_FOoH;N
80FN_k:0RR0FkR8#0_oDFH
O;#:FRR0FkR8#0_oDFH2OR;-

-0RN0LsHkR0C8DCON0sNHRFMVRFs#oHMD#CRFOksCCR8#MHoICNs
RRRRRRRR0N0skHL0#CR$LM_k0HDH8M_kRR:#H0sM
o;RRRRRRRRNs00H0LkC$R#Mk_LHHD0Mk_8RRFV7LW_OR_g:MRC0$H0RRH#"NIC	
";
M
C8WR7__LOg
;
NEsOHO0C0CksRDs0RRFV7LW_OR_gH
#
-N-R0H0sLCk0RO8CDNNs0MHFRsVFRM#HoRDC#sFkO8CRCo#HMsINCNR
0H0sLCk0RM#$_HLkDM0H_R8k:0R#soHM;0
N0LsHkR0C#_$MLDkH0_HM8FkRV0RsDRR:NEsOHO0C0CksRRH#"NIC	
";R-
-RswFRM#HoRDC#sFkO7CRWN,RsHOE00COkRsC#kEFDL8RCkR8l
l$Ns00H0LkC$R#MD_LN_O	LRFG:FRLFNDCMN;
0H0sLCk0RM#$_NLDOL	_FFGRV0RsDRR:NEsOHO0C0CksRRH#0Csk;


LHCoMM
C80RsD
;
-----------------------------------------------------------------------------
-

LDHs$NsR Q  W,7q;) 
Ck#R Q  03#8F_Do_HO4c4n3DND;#
kCWR7q3) 7wW_F8kMNF0HMF_OlNb_sEH03DND;C

M00H$WR7__LO4HjR#F
bs50RO0Nbk_sCORD	:MRHR8#0_oDFH
O;kNb80OC_D:	RRRHM#_08DHFoOO;
Nkb0sCC_MRR:H#MR0D8_FOoH;b
k8CN0_RCM:MRHR8#0_oDFH
O;#VEH0s_8RH:RM0R#8F_Do;HO
8lFCRR:H#MR0D8_FOoH;H
#RH:RM0R#8F_Do;HO
MbH_bHMk:0RRRHM#_08DHFoOF;
kk0b0N_80:NRRRHM#_08DHFoO8;
N_0NFRk0:kRF00R#8F_Do;HO
R#F:kRF00R#8F_DoRHO2
;
-N-R0H0sLCk0RO8CDNNs0MHFRsVFRM#HoRDC#sFkO8CRCo#HMsINCR
RRRRRR0RN0LsHkR0C#_$MLDkH0_HM8:kRRs#0H;Mo
RRRRRRRR0N0skHL0#CR$LM_k0HDH8M_kVRFR_7WL4O_jRR:CHM00H$R#IR"C"N	;


CRM87LW_Oj_4;N

sHOE00COkRsCsR0DF7VRWO_L_R4jH-#
-0RN0LsHkR0C8DCON0sNHRFMVRFs#oHMD#CRFOksCCR8#MHoICNsR0
N0LsHkR0C#_$MLDkH0_HM8:kRRs#0H;Mo
0N0skHL0#CR$LM_k0HDH8M_kVRFRDs0RN:RsHOE00COkRsCH"#RI	CN"R;

R--wRFs#oHMD#CRFOksCWR7,sRNO0EHCkO0s#CREDFk8CRLRl8klN$
0H0sLCk0RM#$_NLDOL	_F:GRRFLFDMCN;0
N0LsHkR0C#_$MLODN	F_LGVRFRDs0RN:RsHOE00COkRsCH0#Rs;kC
C
Lo
HM
8CMRDs0;-

-----------------------------------------------------------------------------


DsHLNRs$Q   ,q7W)7 ,W;jn
Ck#R Q  03#8F_Do_HO4c4n3DND;#
kCWR7q3) 7NWbOo	NCN#3D
D;kR#C7)Wq W37_kwFM08NH_FMN0sHED3NDk;
#7CRW q)3_7WwMFk8HN0FOM_F_lbN0sHED3ND
;
CHM007$RW#_N$HlVV#F_.V_#R
H#oCCMsRHO508NNM_H_8IH0:ERRaQh )t RR:=4
n;8NN0_0Fk_8IH0:ERRaQh )t RR:=U8;
CEb0RQ:Rhta  :)R=nR4;k
b#NE_CP_DDRR:Q hatR ):.=R;k
b#NE_VP_DDRR:Q hatR ):.=R;F
bbC_N_DDPRQ:Rhta  :)R=;R.
bbF__NVDRPD:hRQa  t)=R:R
.;C_sslCF8RQ:Rhta  :)R=;Rj
#bkE$_#M:ORRaQh )t RR:=.b;
F#b_$RMO:hRQa  t)=R:R
.;s_#0lCF8RQ:Rhta  :)R=;R4
0L$Cs_F8RCs:hRQa  t)=R:R2jR;F
bs50RO_D	bEk#RH:RM0R#8F_Do;HO
	OD_bbFRH:RM0R#8F_Do;HO
0s#_:MRRRHM#_08DHFoOb;
k_#Es_CJMRR:H#MR0D8_FOoH;D
Vk_#EMRR:H#MR0D8_FOoH;F
bbC_sJR_M:MRHR8#0_oDFH
O;8NN0_RHM:MRHR8#0_oDFHPO_CFO0sN580HN_MH_I8-0E4FR8IFM0R;j2
#bkEl_CbR0$:kRF00R#8F_Do;HO
#bkEC_NRF:Rk#0R0D8_FOoH;k
b#EE_VRR:FRk0#_08DHFoOb;
k_#EN:VRR0FkR8#0_oDFH
O;bEk#_DVkDRR:FRk0#_08DHFoOs;
NVl_kRDD:kRF00R#8F_Do;HO
sbN08_IRF:Rk#0R0D8_FOoH;k
b#CE_sssFRF:Rk#0R0D8_FOoH;F
bbl_CbR0$:kRF00R#8F_Do;HO
bbF_RNC:kRF00R#8F_Do;HO
bbF_REV:kRF00R#8F_Do;HO
bbF_RNV:kRF00R#8F_Do;HO
bbF_DVkDRR:FRk0#_08DHFoOb;
FCb_sssFRF:Rk#0R0D8_FOoH;N
80FN_k:0RR0FkR8#0_oDFHPO_CFO0sN580FN_kI0_HE80-84RF0IMF2Rj

2;-N-R0H0sLCk0RO8CDNNs0MHFRsVFRM#HoRDC#sFkO8CRCo#HMsINCR
RRRRRR0RN0LsHkR0C#_$MLDkH0_HM8:kRRs#0H;Mo
RRRRRRRR0N0skHL0#CR$LM_k0HDH8M_kVRFR_7WNl#$VFHV__#.#:VRR0CMHR0$H"#RI	CN"C;
M78RW#_N$HlVV#F_.V_#;N

sHOE00COkRsCsR0DF7VRW#_N$HlVV#F_.V_#R
H#-N-R0H0sLCk0RO8CDNNs0MHFRsVFRM#HoRDC#sFkO8CRCo#HMsINCNR
0H0sLCk0RM#$_HLkDM0H_R8k:0R#soHM;0
N0LsHkR0C#_$MLDkH0_HM8FkRV0RsDRR:NEsOHO0C0CksRRH#"NIC	
";
R--wRFs#oHMD#CRFOksCWR7,sRNO0EHCkO0s#CREDFk8CRLRl8klN$
0H0sLCk0RM#$_NLDOL	_F:GRRFLFDMCN;0
N0LsHkR0C#_$MLODN	F_LGVRFRDs0RN:RsHOE00COkRsCH0#Rs;kC
oLCH
M
CRM8s;0D
-
-------------------------------------------------------------------------------------
D

HNLssQ$R ,  7)Wq W,7j
d;kR#CQ   38#0_oDFH4O_43ncN;DD
Ck#Rq7W)7 3WObN	CNo#D3NDk;
#7CRW q)3_7WwMFk8HN0FNM_sEH03DND;#
kCWR7q3) 7wW_F8kMNF0HMF_OlNb_sEH03DND;C

M00H$WR7_$N#lVVHFDO0__#.#HVR#C
oMHCsO
R58NN0__HMI0H8ERR:Q hatR ):c=R;N
80FN_kI0_HE80RQ:Rhta  :)R=nR4;C
8bR0E:hRQa  t)=R:R
U;bEk#__NCDRPD:hRQa  t)=R:R
.;bEk#__NVDRPD:hRQa  t)=R:R
.;b_FbNDC_P:DRRaQh )t RR:=.b;
FNb_VP_DDRR:Q hatR ):.=R;s
CsF_l8:CRRaQh )t RR:=jb;
k_#E#O$MRQ:Rhta  :)R=;R4
bbF_M#$ORR:Q hatR ):4=R;#
s0F_l8:CRRaQh )t RR:=4L;
$_0CFCs8sRR:Q hatR ):j=R

2;b0FsRO5
Db	_kR#E:MRHR8#0_oDFH
O;O_D	bRFb:MRHR8#0_oDFH
O;s_#0MRR:H#MR0D8_FOoH;k
b#sE_CMJ_RH:RM0R#8F_Do;HO
kVD#ME_RH:RM0R#8F_Do;HO
bbF_JsC_:MRRRHM#_08DHFoO8;
N_0NH:MRRRHM#_08DHFoOC_POs0F508NNM_H_8IH04E-RI8FMR0Fj
2;s88_NR0N:MRHR8#0_oDFHPO_CFO0sN5lGkHllN580HN_MH_I8,0E
08NNk_F0H_I820E-84RF0IMF2Rj;C
I_:MRR0FkR8#0_oDFH
O;bEk#_bCl0:$RR0FkR8#0_oDFH
O;bEk#_RNC:kRF00R#8F_Do;HO
#bkEV_ERF:Rk#0R0D8_FOoH;k
b#NE_VRR:FRk0#_08DHFoOb;
k_#EVDkDRF:Rk#0R0D8_FOoH;N
slk_VD:DRR0FkR8#0_oDFH
O;b0Ns_RI8:kRF00R#8F_Do;HO
#bkEs_CsRFs:kRF00R#8F_Do;HO
bbF_bCl0:$RR0FkR8#0_oDFH
O;b_FbN:CRR0FkR8#0_oDFH
O;b_FbE:VRR0FkR8#0_oDFH
O;b_FbN:VRR0FkR8#0_oDFH
O;b_FbVDkDRF:Rk#0R0D8_FOoH;F
bbs_CsRFs:kRF00R#8F_Do;HO
_Is8NN0RF:Rk#0R0D8_FOoH_OPC05FslHNGl5kl8NN0__HMI0H8E8,
N_0NF_k0I0H8E42-RI8FMR0Fj
2;INs_8R8s:kRF00R#8F_Do_HOP0COFLs5HI0_HE805b8C0-E24FR8IFM0R;j2
_s8Ns88RF:Rk#0R0D8_FOoH_OPC05FsL_H0I0H8EC58b20E-84RF0IMF2Rj;N
80FN_k:0RR0FkR8#0_oDFHPO_CFO0sN580FN_kI0_HE80-84RF0IMF2Rj

2;-N-R0H0sLCk0RO8CDNNs0MHFRsVFRM#HoRDC#sFkO8CRCo#HMsINCR
RRRRRR0RN0LsHkR0C#_$MLDkH0_HM8:kRRs#0H;Mo
RRRRRRRR0N0skHL0#CR$LM_k0HDH8M_kVRFR_7WNl#$VFHVO_0D##._VRR:CHM00H$R#IR"C"N	;M
C8WR7_$N#lVVHFDO0__#.#
V;
ONsECH0Os0kC0RsDFRRVWR7_$N#lVVHFDO0__#.#HVR#-

-0RN0LsHkR0C8DCON0sNHRFMVRFs#oHMD#CRFOksCCR8#MHoICNsR0
N0LsHkR0C#_$MLDkH0_HM8:kRRs#0H;Mo
0N0skHL0#CR$LM_k0HDH8M_kVRFRDs0RN:RsHOE00COkRsCH"#RI	CN"
;
-w-RF#sRHDMoCFR#kCsOR,7WRONsECH0Os0kCER#F8kDRRLC8lkl$0
N0LsHkR0C#_$MLODN	F_LGRR:LDFFC;NM
0N0skHL0#CR$LM_D	NO_GLFRRFVsR0D:sRNO0EHCkO0sHCR#sR0k
C;LHCoMC

Ms8R0
D;
---------------------------------------------------------------------------------

-FRBlMbFCRM07#W_J
s0-B-RFNM0HRM#8lkl$sRNO0EHCkO0s
C
DsHLNRs$Q   ,WR7q;) 
Ck#R Q  03#8F_Do_HO4c4n3DND;#
kCWR7q3) 7NWbOo	NCN#3D
D;kR#C7)Wq W37_kwFM08NH_FMObFl_HNs0NE3D
D;
0CMHR0$7#W_JRs0H
#
oCCMsRHO58IH0:ERR#bFHP0HC=R:R;d.
_0OlCF8RM:RNs0kN:DR=2R4;b

FRs05:NRRRHM#_08DHFoOC_POs0F58IH04E-RI8FMR0Fj
2;s0FFRF:Rk#0R0D8_FOoH_OPC05Fs58IH04E+2-/.4FR8IFM0R2j2;-

-0RN0LsHkR0C8DCON0sNHRFMVRFs#oHMD#CRFOksCCR8#MHoICNs
RRRRRRRR0N0skHL0#CR$LM_k0HDH8M_kRR:#H0sM
o;RRRRRRRRNs00H0LkC$R#Mk_LHHD0Mk_8RRFV7#W_JRs0:MRC0$H0RRH#"NIC	
";CRM87#W_J;s0
s
NO0EHCkO0ssCR0FDRVWR7_s#J0#RH
-
-R0N0skHL08CRCNODsHN0FVMRF#sRHDMoCFR#kCsOR#8CHIoMNRsC
0N0skHL0#CR$LM_k0HDH8M_kRR:#H0sM
o;Ns00H0LkC$R#Mk_LHHD0Mk_8RRFVsR0D:sRNO0EHCkO0sHCR#IR"C"N	;-

-FRwsHR#MCoDRk#FsROC7RW,NEsOHO0C0CksRF#EkRD8L8CRk$ll
0N0skHL0#CR$LM_D	NO_GLFRL:RFCFDN
M;Ns00H0LkC$R#MD_LN_O	LRFGFsVR0:DRRONsECH0Os0kC#RHRk0sCL;
CMoH
M
C80RsD
;

-----------------------------------------------------------------------------------------------------
-
R--aDH0CRRRRRRR:WR7_P8H_J#C
R--7HC#oRMRRRRR:WR7_P8H
R--qEk0FRsRRRRR:CR1DlPNR/)RRs]NHR#Ev
Ri-B-RFNlbMR$RR:RRRM1$bODHHR0$10FVICNsR8QMHuNRPR03p308

---------------------------------------------------------------------------------------------------
---7-RCs#OHHb0F:MRR_7W8_HP#RCJHN#RRJ#Ck0CMHRND8HHP8RCs8HC#o8MCRsVFRIDFRCNsNs,NC0N-HRlC08sNCV-FVF,Rs-R
-HREoVERskCJC$MORl5#NRDDOD$OCHR0lRC2NDbbH0ONH#FM3WR7_P8H_J#CRRH#NHMRMo0CC8sRH8PHCIsRHR0ELEF0
R--J0kFH0CMR8NMRlsCN8HMCFsRkk0b0R#3

---------------------------------------------------------------------------------------------------
--SH
DLssN$ RQ 8 ,ICNs;#
kC RQ # 30D8_FOoH_n44cD3NDk;
#HCRC3CC#_08DHFoOM_k#MHoCN83D
D;kR#CHCCC38#0_oDFHNO_sEH03DND;-
-kR#CI	Fs3P8H_J#C_ObN	D3NDk;
#8CRICNs3b7WNNO	o3C#N;DD
Ck#RN8Is7C3WF_wkNM80MHF_lOFbs_NH30EN;DD
C

M00H$WR7_P8H_J#CR
H#SMoCCOsH5S
SNH_I8S0ERm:u1QQae: S=;RU
LSS_8IH0RES:1umQeaQ =S:R
c;SOS0_8lFC:SRQ hatS ):j=R;S
SM_klOR$ORh:Qa  t):RR=;Rd
sSS#l0_FR8C:aQh )t R=R:R
j;SMSHb_k0lCF8Rh:Qa  t)=R:R
4;SkSF00bk_8lFCQR:hta  :)R=;R4
CSSN$sD_N#0s:0RQ hatR ):j=R
2SS;b
SF5s0RSR
S	ODS:SSRRHM#_08DHFoOS;
S0s#_SMRSH:RM0R#8F_Do;HO
ESSFSD8SH:RM0R#8F_Do;HO
#SS00NsSRS:H#MR0D8_FOoH;S
SNSRSSH:RM0R#8F_Do_HOP0COFNs5_8IH04E-RI8FMR0Fj
2;SRSLS:SSRRHM#_08DHFoOC_POs0F5IL_HE80-84RF0IMF2Rj;S
SObFlDCC0SF:Rk#0R0D8_FOoH;SR
SP8HH_8CLj$_SF:Rk#0R0D8_FOoH;S
SJ0kFH0CMSF:Rk#0R0D8_FOoH_OPC05FsNH_I8-0E4FR8IFM0R;j2
sSSCHlNMs8CSF:Rk#0R0D8_FOoH_OPC05FsLH_I8-0E4FR8IFM0R
j2S;S2
-
-R0N0skHL08CRCNODsHN0FVMRF#sRHDMoCFR#kCsOR#8CHIoMN
sCRRRRRRRRNs00H0LkC$R#Mk_LHHD0Mk_8R#:R0MsHoR;
RRRRRNRR0H0sLCk0RM#$_HLkDM0H_R8kF7VRWH_8PC_#JRR:CHM00H$R#IR"C"N	;C

M78RWH_8PC_#J
;
NEsOHO0C0CksRDs0RRFV78W_H#P_CHJR#
R
-N-R0H0sLCk0RO8CDNNs0MHFRsVFRM#HoRDC#sFkO8CRCo#HMsINCNR
0H0sLCk0RM#$_HLkDM0H_R8k:0R#soHM;0
N0LsHkR0C#_$MLDkH0_HM8FkRV0RsDRR:NEsOHO0C0CksRRH#"NIC	
";
R--wRFs#oHMD#CRFOksCWR7,sRNO0EHCkO0s#CREDFk8CRLRl8klN$
0H0sLCk0RM#$_NLDOL	_F:GRRFLFDMCN;0
N0LsHkR0C#_$MLODN	F_LGVRFRDs0RN:RsHOE00COkRsCH0#Rs;kC
C
Lo
HM
CS
Ms8R0
D;

SS
-
-_________________________________________________________________________
__---
-FSv8HHVCL8R$SR:)QqeRDYCDbNbN-
-S07NCSR:SbSqsRHD.Rc,.djj
S--7OC#s0HbHRFM:ESaCsRFHMoHNODRFR8CIRN#VOkM0MHFN$DDROHMFCssOV0RF#sRHCoM8-R
-SSSSbSFC0sNH#FM3aRRECCRsssFRRH#VCHG8FRMIHRI00ERERH#MRCIOCF83-
-
_--_________________________________________________________________________
_

LDHs$NsR Q  I,8N;sC
Ck#R Q  03#8F_Do_HO4c4n3DND;#
kCCRHC#C30D8_FOoH_#kMHCoM8D3NDk;
#HCRC3CC#_08DHFoOs_NH30EN;DD
Ck#RN8Is7C3WObN	CNo#D3NDk;
#8CRICNs3_7WwMFk8HN0FOM_F_lbN0sHED3ND
;
CHM007$RWH_lMGlNR
H#SMoCCOsH5S
SS8IH0RERRRRR:qRhaqz)pR:=dS;
SkSMlM_Hb#k0Rh:Rq)azq=p:RSg
RRRRR2RR;b
SF5s0
NSSRRSRSH:RM#RS0D8_FOoH_OPC05Fs58IH0*ERRlMk_bHMk20#-84RF0IMF2Rj;S
S0ROSRRS:HSMR#_08DHFoOS;
SMlH_GlNRRR:HSMR#_08DHFoOS;
SDPNk:CSR0FkR#RR0D8_FOoH_OPC05FsR8IH04E-RI8FMR0Fj
2;SMSH8SCG:kRF00S#8F_Do_HOP0COFRs5ODCHD.FoRM5RkHl_M0bk#-R24FR8IFM0R
j2S;S2
-
-R0N0skHL08CRCNODsHN0FVMRF#sRHDMoCFR#kCsOR#8CHIoMN
sCRRRRRRRRNs00H0LkC$R#Mk_LHHD0Mk_8R#:R0MsHoR;
RRRRRNRR0H0sLCk0RM#$_HLkDM0H_R8kF7VRWH_lMGlNRC:RM00H$#RHRC"IN;	"
M
C8WR7_MlHlRNG;



ONsECH0Os0kC0RsDVRFR_7WllHMNRGRH
#
-N-R0H0sLCk0RO8CDNNs0MHFRsVFRM#HoRDC#sFkO8CRCo#HMsINCNR
0H0sLCk0RM#$_HLkDM0H_R8k:0R#soHM;0
N0LsHkR0C#_$MLDkH0_HM8FkRV0RsDRR:NEsOHO0C0CksRRH#"NIC	
";
R--wRFs#oHMD#CRFOksCWR7,sRNO0EHCkO0s#CREDFk8CRLRl8klN$
0H0sLCk0RM#$_NLDOL	_F:GRRFLFDMCN;0
N0LsHkR0C#_$MLODN	F_LGVRFRDs0RN:RsHOE00COkRsCH0#Rs;kC
L

CMoH
C

Ms8R0
D;
-
----------------------------------------------------------------------------------------------------
--
-R0aHDRCRRRRRR7:RWH_8P-
-R#7CHRoMRRRRR7:RWH_8P-
-R0qkERFsRRRRR1:RCNDPlRR)/NR]sEH#RivR
R--BbFlNRM$RRRR:$R1MHbDO$H0RV1F0sINCMRQ8RHNu3P0R8p03-
-
---------------------------------------------------------------------------------------------------
R--7OC#s0HbHRFM:WR7_P8HRRH#NFROlMLHNF0HMRNDHCM0oRCs8HHP8RCsIEH0S0LFEkRJFC0HMN0RMs8RCHlNMs8CR0Fkb#k03-R
-ERaHO#RFFlbM0CMRP8HH#8CRC0ERP8HHM8C8N,R,$RLRC0ERP8HHs#F,,RLRR0Fb8sFkROC0RECJ0kFH0CMR8NMRlsCN8HMC
s3-m-RbF0HMDND$0,REsCRCHlNMs8CR0FkbRk0ObFlk#0CRC0ER8lFk#Dk3-
-
R--aREC#MHoRRFV0RECsNClHCM8s#RHRC0ERo#HMVRFRC0ERHqRM0bk3-
-RCaERo#HMVRFRC0ER8lFk#DkRRH#0REC#MHoRRFV0RECAMRHb3k0
---------------------------------------------------------------------------------------------------


SDsHLNRs$Q   ;#
kC RQ # 30D8_FOoH_n44cD3NDk;
#HCRC3CC#_08DHFoOM_k#MHoCN83D
D;kR#CHCCC38#0_oDFHNO_sEH03DND;C

M00H$WR7_P8HR
H#SMoCCOsH5S
SNH_I8S0ERm:u1QQae: S=;4c
LSS_8IH0RES:1umQeaQ =S:gS;
S_0OlCF8ShR:q)azqSpR:;=j
sSSCll_FR8C:ahqzp)qS4:=
2SS;b
SF5s0
NSSRSSS:MRHR8#0_oDFHPO_CFO0s_5NI0H8ER-48MFI0jFR2S;
SSLRSRS:H#MR0D8_FOoH_OPC05FsLH_I8-0E4FR8IFM0R;j2
JSSkHF0CSM0:kRF00R#8F_Do_HOP0COFNs5_8IH04E-RI8FMR0Fj
2;SCSslMNH8SCs:kRF00R#8F_Do_HOP0COFLs5_8IH04E-RI8FMR0Fj
2;SHS8PCH8__L$jRS:FRk0#_08DHFoOS
S2
;
-N-R0H0sLCk0RO8CDNNs0MHFRsVFRM#HoRDC#sFkO8CRCo#HMsINCR
RRRRRR0RN0LsHkR0C#_$MLDkH0_HM8:kRRs#0H;Mo
RRRRRRRR0N0skHL0#CR$LM_k0HDH8M_kVRFR_7W8RHP:MRC0$H0RRH#"NIC	
";
8CMR_7W8RHP;N

sHOE00COkRsCsR0DF7VRWH_8P#RHR-

-0RN0LsHkR0C8DCON0sNHRFMVRFs#oHMD#CRFOksCCR8#MHoICNsR0
N0LsHkR0C#_$MLDkH0_HM8:kRRs#0H;Mo
0N0skHL0#CR$LM_k0HDH8M_kVRFRDs0RN:RsHOE00COkRsCH"#RI	CN"
;
-w-RF#sRHDMoCFR#kCsOR,7WRONsECH0Os0kCER#F8kDRRLC8lkl$0
N0LsHkR0C#_$MLODN	F_LGRR:LDFFC;NM
0N0skHL0#CR$LM_D	NO_GLFRRFVsR0D:sRNO0EHCkO0sHCR#sR0k
C;
oLCH
M

8CMRDs0;



=--=====================================-
-RaR)pFRO8VCRFvsRz_pa7-X
-====================================
==
DS
HNLssQ$R ;  
Ck#R Q  03#8F_Do_HO4c4n3DND;#
kC RQ # 30D8_FOoH_#kMHCoM8D3ND
;
CHM007$RWk_lD80_G#RH
CSoMHCsORR5
ISSHE80R:SRRahqzp)qRR:=cS;
RRRRRSRRbI4_HE80Rh:Rq)azq:pR=RR.
2SS;b
SFRs05S
SNRRRRRRR:MRHR#RR0D8_FOoH_OPC05FsI0H8ER-48MFI0jFR2S;
SRLRRRRRRH:RMRRR#_08DHFoOC_POs0F58IH04E-RI8FMR0Fj
2;SOS0RRRRRRR:HRMRR8#0_oDFH
O;SbS8DRGRRRR:HRMRR8#0_oDFH
O;SsSbFO8k0RR:FRk0R8#0_oDFHPO_CFO0s*5.I0H8ER-48MFI0jFR22
S;-
-R0N0skHL08CRCNODsHN0FVMRF#sRHDMoCFR#kCsOR#8CHIoMN
sCRRRRRRRRNs00H0LkC$R#Mk_LHHD0Mk_8R#:R0MsHoR;
RRRRRNRR0H0sLCk0RM#$_HLkDM0H_R8kF7VRWk_lD80_GRR:CHM00H$R#IR"C"N	;C

M78RWk_lD80_G
;
NEsOHO0C0CksRDs0RRFV7lW_k_D08HGR#
R
-N-R0H0sLCk0RO8CDNNs0MHFRsVFRM#HoRDC#sFkO8CRCo#HMsINCNR
0H0sLCk0RM#$_HLkDM0H_R8k:0R#soHM;0
N0LsHkR0C#_$MLDkH0_HM8FkRV0RsDRR:NEsOHO0C0CksRRH#"NIC	
";
R--wRFs#oHMD#CRFOksCWR7,sRNO0EHCkO0s#CREDFk8CRLRl8klN$
0H0sLCk0RM#$_NLDOL	_F:GRRFLFDMCN;0
N0LsHkR0C#_$MLODN	F_LGVRFRDs0RN:RsHOE00COkRsCH0#Rs;kC
L

CMoH
M
C80RsD
;

--------------------------------------------------------------------------------
--
LDHs$NsR Q  k;
#QCR 3  #_08DHFoO4_4nNc3DRD;RkR
#QCR 3  #_08DHFoOM_k#MHoCN83DRD;RC

M00H$WR7_8N8#_kL8HGR#o
SCsMCH5OR
ISSHE80RRRR:NRM0NksD=R:R;cR
bSS4H_I8R0E:NRM0NksD=R:R
.RSRSRR
2;SsbF0
R5SSSNRRRR:MRHR0R#8F_Do_HOP0COFIs5HE80-84RF0IMF2Rj;S
SLRRRRRRR:MRHR0R#8F_Do_HOP0COFIs5HE80-84RF0IMF2Rj;S
SORH4RRRR:MRHR0R#8F_Do;HO
OSSHR.RR:RRRRHMR8#0_oDFH
O;S8SN8L#kRRR:HRMR#_08DHFoOS;
SR0OSRRRRH:RM#RR0D8_FOoH;S
S#RN0SH:RM#RR0D8_FOoH;S
SNRPoSH:RM#RR0D8_FOoH;S
S8GbDRRS:HRMR#_08DHFoOS;
Sl#kRRS:FRk0#_08DHFoOC_POs0F58IH04E-RI8FMR0FjS2;
OSSFS4R:kRF00R#8F_Do;HO
OSSFS.R:kRF00R#8F_Do
HOS;S2
-
-R0N0skHL08CRCNODsHN0FVMRF#sRHDMoCFR#kCsOR#8CHIoMN
sCRRRRRRRRNs00H0LkC$R#Mk_LHHD0Mk_8R#:R0MsHoR;
RRRRRNRR0H0sLCk0RM#$_HLkDM0H_R8kF7VRW8_N8L#k_R8G:MRC0$H0RRH#"NIC	
";
8CMR_7WN#88k8L_G
;
NEsOHO0C0CksRDs0RRFV7NW_8k8#LG_8RRH#
-
-R0N0skHL08CRCNODsHN0FVMRF#sRHDMoCFR#kCsOR#8CHIoMNRsC
0N0skHL0#CR$LM_k0HDH8M_kRR:#H0sM
o;Ns00H0LkC$R#Mk_LHHD0Mk_8RRFVsR0D:sRNO0EHCkO0sHCR#IR"C"N	;-

-FRwsHR#MCoDRk#FsROC7RW,NEsOHO0C0CksRF#EkRD8L8CRk$ll
0N0skHL0#CR$LM_D	NO_GLFRL:RFCFDN
M;Ns00H0LkC$R#MD_LN_O	LRFGFsVR0:DRRONsECH0Os0kC#RHRk0sC
;
SC
Lo
HM
8CMRDs0;-

-------------------------------------------------------------------------------------------------
-----
-HRa0RDCRRRRRRR:7bW_H8bC_OlN
R--7HC#oRMRRRRR:WR7_bbHCl8_N-O
-kRq0sEFRRRRRRR:1NNLsHHosNHP#RNM1-
-RlBFb$NMRRRRR1:R$DMbH0OH$FR1VN0IsQCRMN8HR0uP30Rp8-3
-NR70RCSRRRRRRR:K$kDR,44Rj.jU-
-
---------------------------------------------------------------------------------------------------
LDHs$NsR Q  W,7q;) 
Ck#R Q  03#8F_Do_HO4c4n3DND;#
kCWR7q3) 7wW_F8kMNF0HMF_OlNb3D
D;
0CMHR0$7bW_H8bC_OlNR
H#
MoCCOsHRS5
NH_I8R0E:mRu1QQae: R=;RU
_SLI0H8ERR:uQm1a QeRR:=US;
N_OOI0H8ERR:uQm1a QeRR:=4
n;SR0O:qRhaqz)p=R:R
j;SbbHCC_soRR:hzqa)Rqp:j=R;H
S8H_I8R0E:mRu1QQae: R=;R4
FSM_Rbl:qRhaqz)p=R:RSj
2
;
b0FsRS5
ORD	:MRHR8#0_oDFH
O;S0s#_:MRRRHM#_08DHFoOS;
H0MH_:MRRRHM#_08DHFoOS;
O_DsN_OOMRR:H#MR0D8_FOoH;N
SRH:RM0R#8F_Do_HOP0COFNs5_8IH04E-RI8FMR0Fj
2;S:LRRRHM#_08DHFoOC_POs0F5IL_HE80-84RF0IMF2Rj;N
SO:ORR0FkR8#0_oDFHPO_CFO0sO5NOH_I8-0E4FR8IFM0R;j2
NSDkEMORH:RM0R#8F_Do;HO
NSDkEMO_RH8:MRHR8#0_oDFHPO_CFO0s85H_8IH04E-RI8FMR0Fj
2;SbbHCk_VD:DRR0FkR8#0_oDFH
O;SbbHCP_FVRR:FRk0#_08DHFoOS;
NCOObM0_RH:RM0R#8F_Do;HO
sSNsCHPRF:Rk#0R0D8_FOoH;N
SsPsHC8_HRF:Rk#0R0D8_FOoH_OPC05FsHI8_HE80-84RF0IMF2Rj;b
Sk_#EF_k0MRR:FRk0#_08DHFoOS;
bCHb_MOC#Rk#:kRF00R#8F_Do_HOP0COF.s5RI8FMR0FjS2
2
;
-N-R0H0sLCk0RO8CDNNs0MHFRsVFRM#HoRDC#sFkO8CRCo#HMsINCR
RRRRRR0RN0LsHkR0C#_$MLDkH0_HM8:kRRs#0H;Mo
RRRRRRRR0N0skHL0#CR$LM_k0HDH8M_kVRFR_7WbCHb8N_lORR:CHM00H$R#IR"C"N	;C

M78RWH_bb_C8l;NO
N

sHOE00COkRsCsR0DF7VRWH_bb_C8lRNOH
#
-N-R0H0sLCk0RO8CDNNs0MHFRsVFRM#HoRDC#sFkO8CRCo#HMsINCNR
0H0sLCk0RM#$_HLkDM0H_R8k:0R#soHM;0
N0LsHkR0C#_$MLDkH0_HM8FkRV0RsDRR:NEsOHO0C0CksRRH#"NIC	
";
R--wRFs#oHMD#CRFOksCWR7,sRNO0EHCkO0s#CREDFk8CRLRl8klN$
0H0sLCk0RM#$_NLDOL	_F:GRRFLFDMCN;0
N0LsHkR0C#_$MLODN	F_LGVRFRDs0RN:RsHOE00COkRsCH0#Rs;kC
LS
CMoH
M
C80RsD
;

