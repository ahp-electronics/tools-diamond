library verilog;
use verilog.vl_types.all;
entity cfg_port is
    generic(
        mst_idle        : integer := 0;
        mst_csdly       : integer := 8;
        mst_mcsn        : integer := 1;
        mst_ldly        : integer := 3;
        mst_mrun        : integer := 2;
        mst_mhld        : integer := 6;
        mst_tdly        : integer := 7;
        mst_rcsn        : integer := 5;
        mst_idly        : integer := 4;
        mst_pcsn        : integer := 9;
        mst_pavn        : integer := 11;
        mst_pavd        : integer := 10;
        mst_pdel1       : integer := 14;
        mst_pdel2       : integer := 15;
        mst_poen        : integer := 13;
        mst_pfin        : integer := 12
    );
    port(
        sfdp_en         : in     vl_logic;
        njbse_sign_read : in     vl_logic;
        njbse_sign_cmd  : in     vl_logic;
        njbse_sign_cmd_read: in     vl_logic;
        sign_match      : out    vl_logic;
        preamblePass    : out    vl_logic;
        signatureCheckEvent: out    vl_logic;
        scanen          : in     vl_logic;
        mclk_byp        : in     vl_logic;
        sck_tcv         : in     vl_logic;
        mclk_int        : in     vl_logic;
        intclk          : in     vl_logic;
        smclk           : in     vl_logic;
        njtrx_rst_async : in     vl_logic;
        njtrx_rst_async0: in     vl_logic;
        tdi             : in     vl_logic;
        cclk_in         : in     vl_logic;
        mclk_in         : in     vl_logic;
        scm_si          : in     vl_logic;
        sspi_si         : in     vl_logic;
        sspi_holdn      : in     vl_logic;
        scpu_writen     : in     vl_logic;
        p16_in          : in     vl_logic_vector(15 downto 0);
        ctrl_mfreq_div  : in     vl_logic_vector(5 downto 0);
        ctrl_lsbf       : in     vl_logic;
        ctrl_cpol       : in     vl_logic;
        ctrl_cpha       : in     vl_logic;
        ctrl_mclk_byp   : in     vl_logic;
        ctrl_tx_edge    : in     vl_logic;
        cfg_ctrl0_upd   : in     vl_logic;
        cfg_mstr_start  : in     vl_logic;
        cfg_mstr_stop   : in     vl_logic;
        cfg_mtx_dat     : in     vl_logic_vector(7 downto 0);
        cfg_mcsn_dat    : in     vl_logic_vector(7 downto 0);
        njbse_sstcmd    : in     vl_logic;
        njbse_txcmd     : in     vl_logic;
        njbse_preamble  : in     vl_logic;
        njbse_rxall     : in     vl_logic;
        njbse_bypass    : in     vl_logic;
        tx_setmcpu      : in     vl_logic;
        tx_command      : in     vl_logic;
        tx_operand      : in     vl_logic;
        restart_bse_en  : in     vl_logic;
        rfifo_full      : in     vl_logic;
        wfifo_empty     : in     vl_logic;
        wfifo_out       : in     vl_logic_vector(15 downto 0);
        jburst_en       : in     vl_logic;
        jburst_pause    : in     vl_logic;
        jburst_01       : in     vl_logic;
        jburst_08       : in     vl_logic;
        nj_rcv_rd_cmd   : in     vl_logic;
        njs_halt        : in     vl_logic;
        p_scm           : in     vl_logic;
        p_sspi          : in     vl_logic;
        p_sp8           : in     vl_logic;
        p_sp16          : in     vl_logic;
        p_mspi_slow     : in     vl_logic;
        p_mspi_fast     : in     vl_logic;
        p_mspi_dual     : in     vl_logic;
        p_mspi_quad     : in     vl_logic;
        p_mp8           : in     vl_logic;
        p_mp16          : in     vl_logic;
        p_mp8_quad      : in     vl_logic;
        p_mp16_quad     : in     vl_logic;
        p_sst           : in     vl_logic;
        p_slave_manu    : in     vl_logic;
        i2c_cfg_active  : in     vl_logic;
        i2c_rfifo_we    : in     vl_logic;
        i2c_rfifo_din   : in     vl_logic_vector(7 downto 0);
        wbc_enable      : in     vl_logic;
        wbc_rfifo_we    : in     vl_logic;
        wbc_rfifo_din   : in     vl_logic_vector(7 downto 0);
        mclk_byp_sel    : out    vl_logic_vector(1 downto 0);
        mclk_div_out    : out    vl_logic;
        mclk_en         : out    vl_logic;
        mclk_pol        : out    vl_logic;
        cfg_port_active : out    vl_logic;
        cfg_cfgrst      : out    vl_logic;
        cfg_rfifo_we    : out    vl_logic;
        cfg_rfifo_w16   : out    vl_logic;
        cfg_rfifo_din   : out    vl_logic_vector(15 downto 0);
        cfg_wfifo_re    : out    vl_logic;
        cfg_wfifo_r16   : out    vl_logic;
        preamble_std    : out    vl_logic;
        preamble_enc    : out    vl_logic;
        preamble_std_ext: out    vl_logic;
        preamble_enc_ext: out    vl_logic;
        njm_tr_next     : out    vl_logic;
        njm_tr_done     : out    vl_logic;
        njm_mcpu_done   : out    vl_logic;
        cfg_mstr_busy   : out    vl_logic;
        sspi_so_1st     : out    vl_logic;
        sspi_oe_1st     : out    vl_logic;
        cfg_mclk_o      : out    vl_logic;
        cfg_mclk_oe     : out    vl_logic;
        cfg_mcsn_o      : out    vl_logic_vector(7 downto 0);
        cfg_mcsn_oe     : out    vl_logic_vector(7 downto 0);
        cfg_data_o      : out    vl_logic_vector(15 downto 0);
        cfg_data_oe     : out    vl_logic_vector(15 downto 0);
        cfg_mclk_byp_o  : out    vl_logic;
        cfg_mclk_byp_oe : out    vl_logic;
        cfg_sd_out      : out    vl_logic;
        cfg_busy_o      : out    vl_logic;
        cfg_busy_oe     : out    vl_logic
    );
end cfg_port;
