-- $Header: //synplicity/map202003lat/mappers/cpld/lib/gen_mach/cmp_lt.vhd#1 $
@ER--O_lbD:0RR8lFkRDCoCCMsFN0sHRVDVCRF#sRksbCODFF50DN0CHORbH#v]qB6jjjv
X2DsHLNRs$Q   ;#
kC RQ # 30D8_FOoH_n44cD3ND
;
CHM00B$Rvpu_a#RH
C
oMHCsOH5I8:0ER0HMCsoC:.=4d
2;
sbF0
5
qR,A:MRHR8#0_oDFHPO_CFO0sH5I8-0E4FR8IFM0R;j2
a
pRF:Rk#0R0D8_FOoH
;
2
M
C8vRBua_p;N

sHOE00COkRsCpBe_vpu_aVRFRuBv_RpaH
#
ObFlFMMC0BRBzt_qAR
RRsbF0R5
RRRRRRqjRRRRRRRRRRRRRRRRRRRRRRRRRRRR:HRRMRRRR71a_tpmQ
B;RRRRRjRARRRRRRRRRRRRRRRRRRRRRRRRRRRRRR:RHRMRRaR17m_pt;QB
RRRRBRRQRhRRRRRRRRRRRRRRRRRRRRRRRRRRRR:RRHMR1RRap7_mBtQ;R
RRRRRBamzRRRRRRRRRRRRRRRRRRRRRRRRR:RRRkRF0RRR1_a7pQmtB
2;CRM8ObFlFMMC0
;
ObFlFMMC0BReBR
RRsbF0R5
RRRRRRXRRRRRRRRRRRRRRRRRRRRRRRRRRRRR:FRRkR0RR71a_tpmQ:BR=jR''
2;CRM8ObFlFMMC0
;
ObFlFMMC0hRQeR
RRsbF0R5
RRRRRRQjRRRRRRRRRRRRRRRRRRRRRRRRRRRR:HRRMRRRR71a_tpmQ
B;RRRRRRRmRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR:RFRk0RaR17m_pt2QB;M
C8FROlMbFC;M0
#

HNoMDNROsRs$RRR:#_08DHFoOC_POs0F5HRI8-0E4FR8IFM0R2jR;H
#oDMNRMOF#j0_R#:R0D8_FOoH;L

CMoH
4Sz:BReBmRu)vaRqRu5XO=>F0M#_2jR;z
S.B:RBqz_tuARmR)av5quR=qj>jq52A,RjA=>5,j2RhBQ=F>OM_#0jB,Rm=za>sONsj$52;R2
dSz:FRVsRRHH4MRRR0FI0H8ER-4oCCMsCN0
zSSd4_p:BRBzt_qAmRu)vaRqRu5q>j=q25H,jRA=5>AHR2,B=Qh>sONsH$5-,42RzBmaO=>N$ss5RH22S;
CRM8oCCMsCN0;z
ScQ:RhueRmR)avRqu5=Qj>NROs5s$I0H8E4R-2m,R=a>p2
;
CRM8pBe_vpu_a
;

