library verilog;
use verilog.vl_types.all;
entity config_register is
    port(
        refresh_out     : in     vl_logic;
        prog_128        : in     vl_logic;
        ext_done        : in     vl_logic;
        idcode          : in     vl_logic_vector(31 downto 0);
        clear_finish    : in     vl_logic;
        start           : in     vl_logic;
        operation       : in     vl_logic;
        wakeup_minus    : in     vl_logic;
        exit_abort      : in     vl_logic;
        illegal_rd      : in     vl_logic;
        functional      : in     vl_logic;
        por             : in     vl_logic;
        tlreset         : in     vl_logic;
        tdi             : in     vl_logic;
        shiftir         : in     vl_logic;
        capir           : in     vl_logic;
        upir            : in     vl_logic;
        tck             : in     vl_logic;
        shiftdr         : in     vl_logic;
        updr            : in     vl_logic;
        capdr           : in     vl_logic;
        selbyp_b        : in     vl_logic;
        selbsr          : in     vl_logic;
        asrout_0        : in     vl_logic;
        dsrout_0        : in     vl_logic;
        bsout_0         : in     vl_logic;
        selasr          : in     vl_logic;
        mnfgshift       : in     vl_logic;
        idcode_o        : in     vl_logic;
        ucode_o         : in     vl_logic;
        progucode_o     : in     vl_logic;
        cmd_ld_ucode    : in     vl_logic;
        cmd_rd_ucode    : in     vl_logic;
        progdone_o      : in     vl_logic;
        erasedone_o     : in     vl_logic;
        progsec_o       : in     vl_logic;
        seldsr          : in     vl_logic;
        test_inst       : in     vl_logic;
        xread_dis_o     : in     vl_logic;
        progctrl0_o     : in     vl_logic;
        vfyctrl0_o      : in     vl_logic;
        status_o        : in     vl_logic;
        cmd_prgm_done_r : in     vl_logic;
        cmd_prgm_done_comp: in     vl_logic;
        cmd_prgm_sec    : in     vl_logic;
        cmd_clear_all_r : in     vl_logic;
        cmd_ld_ctrl0    : in     vl_logic;
        cmd_rd_ctrl0    : in     vl_logic;
        not_edit        : in     vl_logic;
        burst_o         : in     vl_logic;
        vfy_crc_o       : in     vl_logic;
        crc_err         : in     vl_logic;
        id_fail_r       : in     vl_logic;
        non_jtag_config : in     vl_logic;
        read_back       : in     vl_logic;
        cmd_bypass      : in     vl_logic;
        cmd_flow_thru   : in     vl_logic;
        program         : in     vl_logic;
        erase_o         : in     vl_logic;
        mux_clk         : in     vl_logic;
        progen_o        : in     vl_logic;
        xread_en_o      : in     vl_logic;
        wakeup          : in     vl_logic;
        cmd_ctrl0_r     : in     vl_logic_vector(31 downto 0);
        cmd_ucode_r     : in     vl_logic_vector(31 downto 0);
        cmd_crc         : in     vl_logic_vector(15 downto 0);
        seler1          : in     vl_logic;
        seler2          : in     vl_logic;
        er1out          : in     vl_logic;
        er2out          : in     vl_logic;
        break_chain     : in     vl_logic;
        jtag_unprogram  : in     vl_logic;
        jtag_functional : in     vl_logic;
        clear_memory    : in     vl_logic;
        selid           : in     vl_logic;
        cmd_bypass_en   : in     vl_logic;
        edit_mod        : in     vl_logic;
        pcm             : in     vl_logic;
        serial          : in     vl_logic;
        wakeup_clk      : in     vl_logic;
        rti             : in     vl_logic;
        spi_sel         : out    vl_logic_vector(2 downto 0);
        refresh_o       : out    vl_logic;
        mclk_en_r       : out    vl_logic;
        mfgen           : out    vl_logic;
        decomp_en       : out    vl_logic;
        auto_clear      : out    vl_logic;
        mck_freq_switch : out    vl_logic;
        jtag_data       : out    vl_logic;
        jtag_addr       : out    vl_logic;
        instruction     : out    vl_logic_vector(7 downto 0);
        tdo_out         : out    vl_logic;
        tdo_en          : out    vl_logic;
        reg_rd_bus      : out    vl_logic_vector(31 downto 0);
        internal_done   : out    vl_logic;
        done_pupb       : out    vl_logic;
        security        : out    vl_logic;
        freq_sel        : out    vl_logic_vector(5 downto 0);
        freq_div        : out    vl_logic_vector(5 downto 0);
        overload        : out    vl_logic_vector(1 downto 0);
        glb_reg_rd      : out    vl_logic;
        nonjtag_cfg_r   : out    vl_logic;
        read_back_r     : out    vl_logic;
        async_rst       : out    vl_logic;
        error           : out    vl_logic;
        done_reg        : out    vl_logic;
        burst_clear     : out    vl_logic;
        wake_period     : out    vl_logic_vector(2 downto 0);
        init            : out    vl_logic;
        init_r          : out    vl_logic;
        tdi_bscan       : out    vl_logic;
        done_pin_low    : out    vl_logic;
        done_pin_override: out    vl_logic;
        test_cntls      : out    vl_logic_vector(55 downto 0)
    );
end config_register;
