library verilog;
use verilog.vl_types.all;
entity invx1v1s is
    port(
        A               : in     vl_logic;
        Z               : out    vl_logic
    );
end invx1v1s;
