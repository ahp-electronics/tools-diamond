--***************************************************************
-- 4-bit up counters with synchronous clear, asynchronous preset, enable, parallel data load, CAI, and CAO.
-- -XiaoQiu ZHOU
--***************************************************************
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.std_logic_unsigned.ALL;
USE ieee.std_logic_arith.ALL;

ENTITY CBUB4 IS 
    PORT (
        D0  : IN std_logic;
        D1  : IN std_logic;
        D2  : IN std_logic;
        D3  : IN std_logic;
        CAI : IN std_logic;
        CLK : IN std_logic;
        SD  : IN std_logic;
        LD  : IN std_logic;
        EN  : IN std_logic;
        CS  : IN std_logic;
        Q0  : OUT std_logic;
        Q1  : OUT std_logic;
        Q2  : OUT std_logic;
        Q3  : OUT std_logic;
        CAO : OUT std_logic
    );
END CBUB4;

ARCHITECTURE lattice_behav OF CBUB4 IS
    SIGNAL Q_i  : std_logic_vector(3 downto 0);
BEGIN

PROCESS (CLK, SD, LD, D0, D1, D2, D3, EN, CS, CAI)
BEGIN
  IF (SD = '1') THEN
    Q_i <= "1111";    
  ELSIF rising_edge(CLK) THEN
    IF (CS = '1') THEN
      Q_i <= "0000";
    ELSIF (LD = '1') THEN
      Q_i <= D3&D2&D1&D0;	
    ELSIF (CAI = '1' AND EN = '1') THEN
      Q_i <= Q_i + 1;
	  END IF;  
  END IF;
end process;

Q0 <= Q_i(0);
Q1 <= Q_i(1);
Q2 <= Q_i(2);
Q3 <= Q_i(3);
CAO <= CAI AND EN AND Q_i(0) AND Q_i(1) AND Q_i(2) AND Q_i(3);

END lattice_behav;
