--$Header: //synplicity/map202003lat/designware/dw02.vhd#1 $
@E---------------------------------------------------------------------------------------------------

---w-RHRDCRRRRR:RRRj8I.E3P8-
-R#7CHRoMRRRRRB:RFNM0HRM#.LdRNO#HR#7CHWoMNRsCObFlFMMC0
#R-B-RFNlbMR$RR:RRRM1$bODHHR0$Q3MO
R--7CN0RRRRRRRR:kRqo6R.,jR.j-U
-kRq0sEFRRRRRRR:1PCDN)lR
R--e#CsHRFMRRRR:3Rd4-
-
---------------------------------------------------------------------------------------------------
H
DLssN$ RQ 7 ,W q),j7W.k;
#QCR 3  #_08DHFoO4_4nNc3D
D;kR#C7)Wq W37b	NON#oC3DND;#
kCWR7j7.3W_j.ObFlFMMC0N#3D
D;
0CMHR0$7.Wj_M#HR
H#oCCMsRHO5_RqI0H8ERR:Q hatR ):4=Rn#;
HIM_HE80RQ:Rhta  :)R=.RdR
2;b0FsRq5RRH:RM0R#8F_Do_HOP0COFqs5_8IH04E-RI8FMR0Fj
2;1RQh:kRF00R#8F_Do_HOP0COF#s5HIM_HE80-84RF0IMF2RjR
2;
-
-R0N0skHL08CRCNODsHN0FVMRF#sRHDMoCFR#kCsOR#8CHIoMN
sCRRRRRRRRNs00H0LkC$R#Mk_LHHD0Mk_8R#:R0MsHoR;
RRRRRNRR0H0sLCk0RM#$_HLkDM0H_R8kF7VRW_j.#RHM:MRC0$H0RRH#"NIC	
";
8CMRj7W.H_#M
;
NEsOHO0C0CksRDs0RRFV7.Wj_M#HR
H#
-R-R0N0skHL08CRCNODsHN0FVMRF#sRHDMoCFR#kCsOR#8CHIoMNRsC
RRRRRRRR0N0skHL0#CR$LM_k0HDH8M_kRR:#H0sM
o;RRRRRRRRNs00H0LkC$R#Mk_LHHD0Mk_8RRFVsR0D:sRNO0EHCkO0sHCR#IR"C"N	;-

-FRwsHR#MCoDRk#FsROC7RW,NEsOHO0C0CksRF#EkRD8L8CRk$ll
0SN0LsHkR0C#_$MLODN	F_LGRR:LDFFC;NM
0SN0LsHkR0C#_$MLODN	F_LGVRFRDs0RN:RsHOE00COkRsCH0#Rs;kC
oLCH
M
CRM8s;0D
-
------------------------------------------------------------------D

HNLssQ$R ,  7)Wq W,7j
.;kR#CQ   38#0_oDFH4O_43ncN;DD
Ck#Rq7W)7 3WObN	CNo#D3NDk;
#7CRW3j.7.Wj_lOFbCFMM30#N;DD
M
C0$H0Rj7W.H_#M#OFR
H#
MoCCOsHRq5R_8IH0:ERRaQh )t RR:=4
n;ICNP_8IH0:ERRaQh )t RR:=d2.R;b

FRs05RRq:MRHR8#0_oDFHPO_CFO0s_5qI0H8ER-48MFI0jFR21;
QBh_m:1RRRHM#_08DHFoOW;
qRe :kRF00R#8F_Do_HOP0COFIs5N_PCI0H8ER-48MFI0jFR2;R2
-
-R0N0skHL08CRCNODsHN0FVMRF#sRHDMoCFR#kCsOR#8CHIoMN
sCRRRRRRRRNs00H0LkC$R#Mk_LHHD0Mk_8R#:R0MsHoR;
RRRRRNRR0H0sLCk0RM#$_HLkDM0H_R8kF7VRW_j.#OHMF:#RR0CMHR0$H"#RI	CN"
;
CRM87.Wj_M#HO;F#
s
NO0EHCkO0ssCR0FDRVWR7j#._HFMO##RH
-
R-0RN0LsHkR0C8DCON0sNHRFMVRFs#oHMD#CRFOksCCR8#MHoICNsRR
RRRRRR0RN0LsHkR0C#_$MLDkH0_HM8:kRRs#0H;Mo
RRRRRRRR0N0skHL0#CR$LM_k0HDH8M_kVRFRDs0RN:RsHOE00COkRsCH"#RI	CN"
;
-w-RF#sRHDMoCFR#kCsOR,7WRONsECH0Os0kCER#F8kDRRLC8lkl$N
S0H0sLCk0RM#$_NLDOL	_F:GRRFLFDMCN;N
S0H0sLCk0RM#$_NLDOL	_FFGRV0RsDRR:NEsOHO0C0CksRRH#0Csk;L

CMoH
8CMRDs0;-

-------------------------------------------------------------------------D

HNLssQ$R ,  7)Wq W,7j
.;kR#CQ   38#0_oDFH4O_43ncN;DD
Ck#Rq7W)7 3WObN	CNo#D3NDk;
#7CRW3j.7.Wj_lOFbCFMM30#N;DD
M
C0$H0Rj7W.F_O##RH
C
oMHCsORR5qH_I8R0E:hRQa  t)=R:R;4n
#OF_8IH0:ERRaQh )t RR:=d2.R;b

FRs05RRq:MRHR8#0_oDFHPO_CFO0s_5qI0H8ER-48MFI0jFR2B;
m:1RR0FkR8#0_oDFHPO_CFO0sF5O#H_I8-0E4FR8IFM0RRj22
;
-N-R0H0sLCk0RO8CDNNs0MHFRsVFRM#HoRDC#sFkO8CRCo#HMsINCR
RRRRRR0RN0LsHkR0C#_$MLDkH0_HM8:kRRs#0H;Mo
RRRRRRRR0N0skHL0#CR$LM_k0HDH8M_kVRFRj7W.F_O#RR:CHM00H$R#IR"C"N	;C

M78RW_j.O;F#
s
NO0EHCkO0ssCR0FDRVWR7jO._FH#R#-
R-0RN0LsHkR0C8DCON0sNHRFMVRFs#oHMD#CRFOksCCR8#MHoICNsRR
RRRRRR0RN0LsHkR0C#_$MLDkH0_HM8:kRRs#0H;Mo
RRRRRRRR0N0skHL0#CR$LM_k0HDH8M_kVRFRDs0RN:RsHOE00COkRsCH"#RI	CN"
;
-w-RF#sRHDMoCFR#kCsOR,7WRONsECH0Os0kCER#F8kDRRLC8lkl$N
S0H0sLCk0RM#$_NLDOL	_F:GRRFLFDMCN;N
S0H0sLCk0RM#$_NLDOL	_FFGRV0RsDRR:NEsOHO0C0CksRRH#0Csk;C
Lo
HM
8CMRDs0;-

-========================================C==M00H$MRN8sRNO0EHCkO0sVCRF8sRI_j.l0kD_#._0CNoR========================D=
HNLssH$RC;CC
Ck#RCHCC03#8F_Do_HO4c4n3DND;#
kCCRHC#C30D8_FOoH_#kMHCoM8D3ND
;
CHM007$RW_j.l0kD_#._0CNoR
H#SMoCCOsH5q
S_8IH0:ERR1umQeaQ 4:=n
R;SIA_HE80Ru:Rma1QQ:e =
4nS
2;b0Fs5q
SR:SSRRHM#_08DHFoOC_POs0F5Iq_HE80-84RF0IMF2Rj;A
SR:SSRRHM#_08DHFoOC_POs0F5IA_HE80-84RF0IMF2Rj;a
SBSRS:MRHR8#0_oDFH
O;SiBpRRS:H#MR0D8_FOoH;u
S)zm7B:aRR0FkR8#0_oDFHPO_CFO0s_5qI0H8E_+AI0H8ER-48MFI0jFR22
S;-
-R0N0skHL08CRCNODsHN0FVMRF#sRHDMoCFR#kCsOR#8CHIoMN
sCRRRRRRRRNs00H0LkC$R#Mk_LHHD0Mk_8R#:R0MsHoR;
RRRRRNRR0H0sLCk0RM#$_HLkDM0H_R8kF7VRW_j.l0kD_#._0CNoRC:RM00H$#RHRC"IN;	"
M
C8WR7jl._k_D0.0_#N;oC
N

sHOE00COkRsCsR0DF7VRW_j.l0kD_#._0CNoR
H#
-R-R0N0skHL08CRCNODsHN0FVMRF#sRHDMoCFR#kCsOR#8CHIoMNRsC
RRRRRRRR0N0skHL0#CR$LM_k0HDH8M_kRR:#H0sM
o;RRRRRRRRNs00H0LkC$R#Mk_LHHD0Mk_8RRFVsR0D:sRNO0EHCkO0sHCR#IR"C"N	;-

-FRwsHR#MCoDRk#FsROC7RW,NEsOHO0C0CksRF#EkRD8L8CRk$ll
0SN0LsHkR0C#_$MLODN	F_LGRR:LDFFC;NM
0SN0LsHkR0C#_$MLODN	F_LGVRFRDs0RN:RsHOE00COkRsCH0#Rs;kC
C
Lo
HM
8CMRDs0;


-=-=========================================CHM00N$RMN8RsHOE00COkRsCVRFs8.Ij_Dlk0__d#o0NC=R======================R==
D

HNLssH$RC;CC
Ck#RCHCC03#8F_Do_HO4c4n3DND;#
kCCRHC#C30D8_FOoH_#kMHCoM8D3ND
;
CHM007$RW_j.l0kD_#d_0CNoR
H#S
SSSMoCCOsH5S
SSIq_HE80Ru:Rma1QQ:e =R4n;S
SSIA_HE80Ru:Rma1QQ:e =
4nS2SS;S
Sb0Fs5S
SSSqRSH:RM0R#8F_Do_HOP0COFqs5_8IH04E-RI8FMR0Fj
2;SASSR:SSRRHM#_08DHFoOC_POs0F5IA_HE80-84RF0IMF2Rj;S
SSRaBSRS:H#MR0D8_FOoH;S
SSiBpRRS:H#MR0D8_FOoH;S
SSmu)7azBRF:Rk#0R0D8_FOoH_OPC05FsqH_I8+0EAH_I8-0E4FR8IFM0R
j2S2SS;-

-0RN0LsHkR0C8DCON0sNHRFMVRFs#oHMD#CRFOksCCR8#MHoICNs
RRRRRRRR0N0skHL0#CR$LM_k0HDH8M_kRR:#H0sM
o;RRRRRRRRNs00H0LkC$R#Mk_LHHD0Mk_8RRFV7.Wj_Dlk0__d#o0NCRR:CHM00H$R#IR"C"N	;C

M78RW_j.l0kD_#d_0CNo;


SsSNO0EHCkO0ssCR0FDRVWR7jl._k_D0d0_#NRoCH
#R
R--Ns00H0LkCCR8OsDNNF0HMFRVsHR#MCoDRk#FsROC8HC#oNMIs
CRRRRRRRRRNs00H0LkC$R#Mk_LHHD0Mk_8R#:R0MsHoR;
RRRRRNRR0H0sLCk0RM#$_HLkDM0H_R8kFsVR0:DRRONsECH0Os0kC#RHRC"IN;	"
-
-RswFRM#HoRDC#sFkO7CRWN,RsHOE00COkRsC#kEFDL8RCkR8l
l$S0N0skHL0#CR$LM_D	NO_GLFRL:RFCFDN
M;S0N0skHL0#CR$LM_D	NO_GLFRRFVsR0D:sRNO0EHCkO0sHCR#sR0k
C;

SSSLS
CMoH
M
C80RsD
;SSRRR
RSRRR
SR
R

=--=========================================0CMHR0$NRM8NEsOHO0C0CksRsVFRj8I.k_lDc0__N#0o=CR========================RD

HNLssH$RC;CC
Ck#RCHCC03#8F_Do_HO4c4n3DND;#
kCCRHC#C30D8_FOoH_#kMHCoM8D3ND
;
SMSC0$H0Rj7W.k_lDc0__N#0oHCR#S
SSMoCCOsHRS5
SqSS_8IH0:ERR0HMCsoCRR:=4
n;SSSSAH_I8R0E:MRH0CCos=R:R
4nSSSSS
2;SbSSFRs05S
SSRSqS:SSRRHM#_08DHFoOC_POs0F5Iq_HE80-84RF0IMF2Rj;S
SSRSAS:SSRRHM#_08DHFoOC_POs0F5IA_HE80-84RF0IMF2Rj;S
SSBSaRRSRR:RSRRHM#_08DHFoOS;
SBSSpSiRSH:RM0R#8F_Do;HO
SSSSmu)7azBRRS:FRk0#_08DHFoOC_POs0F5Iq_HE80+IA_HE80-84RF0IMF2Rj
SSSS
2;
R--Ns00H0LkCCR8OsDNNF0HMFRVsHR#MCoDRk#FsROC8HC#oNMIsRC
RRRRRNRR0H0sLCk0RM#$_HLkDM0H_R8k:0R#soHM;R
RRRRRR0RN0LsHkR0C#_$MLDkH0_HM8FkRVWR7jl._k_D0c0_#NRoC:MRC0$H0RRH#"NIC	
";
CSSM78RW_j.l0kD_#c_0CNo;


SsSNO0EHCkO0ssCR0FDRVWR7jl._k_D0c0_#NRoCH
#
-N-R0H0sLCk0RO8CDNNs0MHFRsVFRM#HoRDC#sFkO8CRCo#HMsINCRR
RRRRRNRR0H0sLCk0RM#$_HLkDM0H_R8k:0R#soHM;R
RRRRRR0RN0LsHkR0C#_$MLDkH0_HM8FkRV0RsDRR:NEsOHO0C0CksRRH#"NIC	
";
R--wRFs#oHMD#CRFOksCWR7,sRNO0EHCkO0s#CREDFk8CRLRl8klS$
Ns00H0LkC$R#MD_LN_O	LRFG:FRLFNDCMS;
Ns00H0LkC$R#MD_LN_O	LRFGFsVR0:DRRONsECH0Os0kC#RHRk0sC
;

oLCH
M

8CMRDs0;R
SR
R
-=-=========================================CHM00N$RMN8RsHOE00COkRsCVRFs8.Ij_Dlk0__6#o0NC=R======================R==
D

HNLssH$RC;CC
Ck#RCHCC03#8F_Do_HO4c4n3DND;#
kCCRHC#C30D8_FOoH_#kMHCoM8D3ND
;
SMSC0$H0Rj7W.k_lD60__N#0oHCR#S
SSMoCCOsHRS5
SqSS_8IH0:ERR0HMCsoCRR:=4
n;SSSSAH_I8R0E:MRH0CCos=R:R
4nSSSSS
2;SbSSFRs05S
SSRSqS:SSRRHM#_08DHFoOC_POs0F5Iq_HE80-84RF0IMF2Rj;S
SSRSAS:SSRRHM#_08DHFoOC_POs0F5IA_HE80-84RF0IMF2Rj;S
SSBSaRRSRR:RSRRHM#_08DHFoOS;
SBSSpSiRSH:RM0R#8F_Do;HO
SSSSmu)7azBRRS:FRk0#_08DHFoOC_POs0F5Iq_HE80+IA_HE80-84RF0IMF2Rj
SSSS
2;
R--Ns00H0LkCCR8OsDNNF0HMFRVsHR#MCoDRk#FsROC8HC#oNMIsRC
RRRRRNRR0H0sLCk0RM#$_HLkDM0H_R8k:0R#soHM;R
RRRRRR0RN0LsHkR0C#_$MLDkH0_HM8FkRVWR7jl._k_D060_#NRoC:MRC0$H0RRH#"NIC	
";
CSSM78RW_j.l0kD_#6_0CNo;


SsSNO0EHCkO0ssCR0FDRVWR7jl._k_D060_#NRoCH
#
-N-R0H0sLCk0RO8CDNNs0MHFRsVFRM#HoRDC#sFkO8CRCo#HMsINCRR
RRRRRNRR0H0sLCk0RM#$_HLkDM0H_R8k:0R#soHM;R
RRRRRR0RN0LsHkR0C#_$MLDkH0_HM8FkRV0RsDRR:NEsOHO0C0CksRRH#"NIC	
";
R--wRFs#oHMD#CRFOksCWR7,sRNO0EHCkO0s#CREDFk8CRLRl8klS$
Ns00H0LkC$R#MD_LN_O	LRFG:FRLFNDCMS;
Ns00H0LkC$R#MD_LN_O	LRFGFsVR0:DRRONsECH0Os0kC#RHRk0sC
;

oLCH
M
S
RRCRM8s;0D
-
-=========================================M=C0$H0R8NMRONsECH0Os0kCFRVsIR8jl._k_D0n0_#NRoC=========================
R

LDHs$NsRCHCCk;
#HCRC3CC#_08DHFoO4_4nNc3D
D;kR#CHCCC38#0_oDFHkO_Mo#HM3C8N;DD
S
SCHM007$RW_j.l0kD_#n_0CNoR
H#SoSSCsMCH5OR
SSSSIq_HE80RH:RMo0CC:sR=nR4;S
SS_SAI0H8ERR:HCM0oRCs:4=RnS
SS2SS;S
SSsbF0
R5SSSSqSRSSH:RM0R#8F_Do_HOP0COFqs5_8IH04E-RI8FMR0Fj
2;SSSSASRSSH:RM0R#8F_Do_HOP0COFAs5_8IH04E-RI8FMR0Fj
2;SSSSaSBRRRRRSH:RM0R#8F_Do;HO
SSSSiBpR:SSRRHM#_08DHFoOS;
SuSS)zm7BSaR:kRF00R#8F_Do_HOP0COFqs5_8IH0AE+_8IH04E-RI8FMR0FjS2
S2SS;-

-0RN0LsHkR0C8DCON0sNHRFMVRFs#oHMD#CRFOksCCR8#MHoICNs
RRRRRRRR0N0skHL0#CR$LM_k0HDH8M_kRR:#H0sM
o;RRRRRRRRNs00H0LkC$R#Mk_LHHD0Mk_8RRFV7.Wj_Dlk0__n#o0NCRR:CHM00H$R#IR"C"N	;S

S8CMRj7W.k_lDn0__N#0o
C;
S
SNEsOHO0C0CksRDs0RRFV7.Wj_Dlk0__n#o0NC#RH
-
-R0N0skHL08CRCNODsHN0FVMRF#sRHDMoCFR#kCsOR#8CHIoMNRsC
RRRRRRRR0N0skHL0#CR$LM_k0HDH8M_kRR:#H0sM
o;RRRRRRRRNs00H0LkC$R#Mk_LHHD0Mk_8RRFVsR0D:sRNO0EHCkO0sHCR#IR"C"N	;-

-FRwsHR#MCoDRk#FsROC7RW,NEsOHO0C0CksRF#EkRD8L8CRk$ll
0SN0LsHkR0C#_$MLODN	F_LGRR:LDFFC;NM
0SN0LsHkR0C#_$MLODN	F_LGVRFRDs0RN:RsHOE00COkRsCH0#Rs;kC
L

CMoH
M
C80RsDR;R
-
----------------------------------------------------------------------
-
DsHLNRs$HCCC;#
kCCRHC#C30D8_FOoH_n44cD3NDk;
#HCRC3CC#_08DHFoOM_k#MHoCN83D
D;kR#CHCCC38#0_oDFHNO_sEH03DND;C

M00H$WR7_k#JNbsCRRH#
CSoMHCsOH5I8R0ERRR:hzqa)Rqp:n=R
RSRRRRRRR2;R
RRSsbF0S5
SRNRRRR:HRMR#_08DHFoOC_POs0F58IH04E-RI8FMR0FjR2;RRRRRRRRSS
S0RORRH:RM#RR0D8_FOoH;
RSSkSF0:jRR0FkR8#0_oDFHPO_CFO0s*5.I0H8ER-48MFI0jFR2S;
S0Fk4RR:FRk0#_08DHFoOC_POs0F5I.*HE80-84RF0IMF2Rj2
;
-N-R0H0sLCk0RO8CDNNs0MHFRsVFRM#HoRDC#sFkO8CRCo#HMsINCR
RRRRRR0RN0LsHkR0C#_$MLDkH0_HM8:kRRs#0H;Mo
RRRRRRRR0N0skHL0#CR$LM_k0HDH8M_kVRFR_7W#NJksRCb:MRC0$H0RRH#"NIC	
";
8CMR_7W#NJks;Cb
s
NO0EHCkO0ssCR0FDRVWR7_k#JNbsCRRH#
-
-R0N0skHL08CRCNODsHN0FVMRF#sRHDMoCFR#kCsOR#8CHIoMNRsC
RRRRRRRR0N0skHL0#CR$LM_k0HDH8M_kRR:#H0sM
o;RRRRRRRRNs00H0LkC$R#Mk_LHHD0Mk_8RRFVsR0D:sRNO0EHCkO0sHCR#IR"C"N	;-

-FRwsHR#MCoDRk#FsROC7RW,NEsOHO0C0CksRF#EkRD8L8CRk$ll
0SN0LsHkR0C#_$MLODN	F_LGRR:LDFFC;NM
0SN0LsHkR0C#_$MLODN	F_LGVRFRDs0RN:RsHOE00COkRsCH0#Rs;kC
L

CMoH
C

Ms8R0
D;
=--=========================================0CMHR0$NRM8NEsOHO0C0CksRsVFRj7W.)_a = R========================
D

HNLssH$RC;CC
Ck#RCHCC03#8F_Do_HO4c4n3DND; 

haaQYWR7j0._sRCCQ
1
RtRR )h Q5BRHkMb0H_I8R0E:hRQa  t)6:=RR;RM_klHkMb0:#RRaQh )t :R=c2R;R
RRRRRR
RmRu)Ra5QzhuaSRSRQ:RhRRR1_a7pQmtB _eB)amRH55M0bk_8IH0ME*kHl_M0bk#42-R7RRmaWhm2Rj;R
RRRRRRmRRz,ajm4zaR:RRRamzRaR17m_pt_QBea Bm5)RHkMb0H_I8-0E4mR7WmhaR2j2;
R
-N-R0H0sLCk0RO8CDNNs0MHFRsVFRM#HoRDC#sFkO8CRCo#HMsINCR
RRRRRR0RN0LsHkR0C#_$MLDkH0_HM8:kRRs#0H;Mo
RRRRRRRR0N0skHL0#CR$LM_k0HDH8M_kVRFRj7W.s_0C:CRR0CMHR0$H"#RI	CN"
;

7 hRj7W.s_0C
C;
)
qBa]Q zBa)s R0FDRVWR7j0._sRCCHR#R
-
-R0N0skHL08CRCNODsHN0FVMRF#sRHDMoCFR#kCsOR#8CHIoMNRsC
RRRRRRRR0N0skHL0#CR$LM_k0HDH8M_kRR:#H0sM
o;RRRRRRRRNs00H0LkC$R#Mk_LHHD0Mk_8RRFVsR0D:sRNO0EHCkO0sHCR#IR"C"N	;-

-FRwsHR#MCoDRk#FsROC7RW,NEsOHO0C0CksRF#EkRD8L8CRk$ll
0SN0LsHkR0C#_$MLODN	F_LGRR:LDFFC;NM
0SN0LsHkR0C#_$MLODN	F_LGVRFRDs0RN:RsHOE00COkRsCH0#Rs;kC
C
LoRHMRS


8CMRDs0;



S--============SMSC0$H0R8NMRONsECH0Os0kCFRVsWR7jv._zupaS=R==========
=

LDHs$NsRCHCCk;
#HCRC3CC#_08DHFoO4_4nNc3D
D;kR#CHCCC38#0_oDFHkO_Mo#HM3C8N;DDS
RRkR#CHCCC38#0_oDFHNO_sEH03DND;C

M00H$WR7jl._kbD0RRH#
CSoMHCsOS5
SIN_HE80R:RRRahqzp)qRR:=nS;
SIL_HE80R:RRRahqzp)qRR:=US;
S0Fk_8IH0:ERRahqzp)qRR:=4SU
SR2;RSR
b0Fs5S
SNRRRRH:RM#RR0D8_FOoH_OPC05FsNH_I8-0E4FR8IFM0R;j2
LSSRRRR:MRHR0R#8F_Do_HOP0COFLs5_8IH04E-RI8FMR0Fj
2;SOS0R:RRRRHMR8#0_oDFHRO;
FSSkR0j:kRF00R#8F_Do_HOP0COFFs5kI0_HE80-84RF0IMF2Rj;S
SF4k0RF:Rk#0R0D8_FOoH_OPC05FsF_k0I0H8ER-48MFI0jFR2S
S2-;
-0RN0LsHkR0C8DCON0sNHRFMVRFs#oHMD#CRFOksCCR8#MHoICNs
RRRRRRRR0N0skHL0#CR$LM_k0HDH8M_kRR:#H0sM
o;RRRRRRRRNs00H0LkC$R#Mk_LHHD0Mk_8RRFV7.Wj_Dlk0:bRR0CMHR0$H"#RI	CN"
;
CRM87.Wj_Dlk0
b;
ONsECH0Os0kC0RsDVRFRj7W.k_lDR0bH
#R
R--Ns00H0LkCCR8OsDNNF0HMFRVsHR#MCoDRk#FsROC8HC#oNMIs
CRRRRRRRRRNs00H0LkC$R#Mk_LHHD0Mk_8R#:R0MsHoR;
RRRRRNRR0H0sLCk0RM#$_HLkDM0H_R8kFsVR0:DRRONsECH0Os0kC#RHRC"IN;	"
-
-RswFRM#HoRDC#sFkO7CRWN,RsHOE00COkRsC#kEFDL8RCkR8l
l$S0N0skHL0#CR$LM_D	NO_GLFRL:RFCFDN
M;S0N0skHL0#CR$LM_D	NO_GLFRRFVsR0D:sRNO0EHCkO0sHCR#sR0k
C;
oLCH
M
CRM8s;0D
-

-========================================C==M00H$MRN8sRNO0EHCkO0sVCRF7sRW_j.b8sF_l#k4=R======================
==DsHLNRs$Q   ;#
kC RQ # 30D8_FOoH_n44cD3NDk;
#HCRC3CC#_08DHFoOM_k#MHoCN83D
D;kR#CHCCC38#0_oDFHNO_sEH03DND;M
C0$H0Rj7W.s_bF#8_kRl4Ho#
CsMCH5OR
qSS_8IH0RERRh:Rq)azq:pR=
d;S_SAI0H8ERRR:qRhaqz)p=R:dS;
Sv1z_8IH0:ERRahqzp)qRc:=
2SS;b
SF5s0
qSSRRS:H#MR0D8_FOoH_OPC05FsqH_I8-0E4FR8IFM0R;j2
ASSRRS:H#MR0D8_FOoH_OPC05FsAH_I8-0E4FR8IFM0R;j2
BSSRRS:H#MR0D8_FOoH_OPC05Fs1_zvI0H8ER-48MFI0jFR2S;
SRaBSH:RM0R#8F_Do;HO
1SSz:vSR0FkR8#0_oDFHPO_CFO0sz51vH_I8-0E4FR8IFM0R
j2SRRRR
2;
R--Ns00H0LkCCR8OsDNNF0HMFRVsHR#MCoDRk#FsROC8HC#oNMIsRC
RRRRRNRR0H0sLCk0RM#$_HLkDM0H_R8k:0R#soHM;R
RRRRRR0RN0LsHkR0C#_$MLDkH0_HM8FkRVWR7jb._s_F8#4klRC:RM00H$#RHRC"IN;	"
M
C8WR7jb._s_F8#4kl;N

sHOE00COkRsCsR0DF7VRW_j.b8sF_l#k4#RH
o#HMRNDb8sFR#:R0D8_FOoH_OPC05FsNH_I8+0ELH_I8-0E4FR8IFM0R;j2SRRR
o#HMRND#MHoLRH0:8#0_oDFH
O;
R--Ns00H0LkCCR8OsDNNF0HMFRVsHR#MCoDRk#FsROC8HC#oNMIs
CRRRRRRRRRNs00H0LkC$R#Mk_LHHD0Mk_8R#:R0MsHoR;
RRRRRNRR0H0sLCk0RM#$_HLkDM0H_R8kFsVR0:DRRONsECH0Os0kC#RHRC"IN;	"
-
-RswFRM#HoRDC#sFkO7CRWN,RsHOE00COkRsC#kEFDL8RCkR8l
l$S0N0skHL0#CR$LM_D	NO_GLFRL:RFCFDN
M;S0N0skHL0#CR$LM_D	NO_GLFRRFVsR0D:sRNO0EHCkO0sHCR#sR0k
C;
C
Lo
HM
8CMRDs0;



-
-=========================================M=C0$H0R8NMRONsECH0Os0kCFRVsWR7j#._k=lR========================
LDHs$NsR Q  k;
#QCR 3  #_08DHFoO4_4nNc3D
D;kR#CHCCC38#0_oDFHkO_Mo#HM3C8N;DD
M
C0$H0Rj7W.k_#l#RH
C
oMHCsOS5
SbHMkI0_HE80Rq:haqz)p=R:cS;
SlMk_bHMkR0#Rq:haqz)p=R:cS
S2S;
b0Fs5S
SQzhuaRS:HRMR#_08DHFoOC_POs0F5bHMkI0_HE80RM*RkHl_M0bk#R-48MFI0jFR2S;
Sv1zR:RSR0FkR8#0_oDFHPO_CFO0sM5Hb_k0I0H8ER-48MFI0jFR2S
S2
;
-N-R0H0sLCk0RO8CDNNs0MHFRsVFRM#HoRDC#sFkO8CRCo#HMsINCR
RRRRRR0RN0LsHkR0C#_$MLDkH0_HM8:kRRs#0H;Mo
RRRRRRRR0N0skHL0#CR$LM_k0HDH8M_kVRFRj7W.k_#lRR:CHM00H$R#IR"C"N	;C

M78RW_j.#;kl
N

sHOE00COkRsCsR0DF7VRW_j.#RklH##
HNoMDkRMlM_Hb#k0_o#HRh:RNs0kN
D;
R--Ns00H0LkCCR8OsDNNF0HMFRVsHR#MCoDRk#FsROC8HC#oNMIs
CRRRRRRRRRNs00H0LkC$R#Mk_LHHD0Mk_8R#:R0MsHoR;
RRRRRNRR0H0sLCk0RM#$_HLkDM0H_R8kFsVR0:DRRONsECH0Os0kC#RHRC"IN;	"
-
-RswFRM#HoRDC#sFkO7CRWN,RsHOE00COkRsC#kEFDL8RCkR8l
l$S0N0skHL0#CR$LM_D	NO_GLFRL:RFCFDN
M;S0N0skHL0#CR$LM_D	NO_GLFRRFVsR0D:sRNO0EHCkO0sHCR#sR0k
C;
oLCHSM

8CMRDs0;


-=-=============S0CMHR0$NRM8NEsOHO0C0CksRsVFRj7W.s_bF#8_k=lS============
H
DLssN$ RQ 
 ;kR#CQ   38#0_oDFH4O_43ncN;DD
Ck#RCHCC03#8F_Do_HOkHM#o8MC3DND;#
kCCRHC#C30D8_FOoH_HNs0NE3D
D;
0CMHR0$7.Wj_Fbs8k_#l#RHRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRS

oCCMsRHO5S
SS_RqI0H8E:RSRahqzp)qRR:=6
R;SRSSAH_I8R0ESh:Rq)azq:pR=RR6;S
SSkRMlM_Hb#k0Su:Rma1QQRe :d=RRS;
S1SRzIv_HE80RRS:hzqa)Rqp:4=R.S
SS
2;SFSbs
05SqSSRRS:H#MR0D8_FOoH_OPC05FsM_klHkMb0*#RRIq_HE80-84RF0IMF2Rj;S
SSSAR:MRHR8#0_oDFHPO_CFO0sk5MlM_Hb#k0RA*R_8IH04E-RI8FMR0Fj
2;SaSSB:RSRRHM#_08DHFoOS;
SzS1vRR:FRk0#_08DHFoOC_POs0F5v1z_8IH04E-RI8FMR0FjS2
SR2;RRRRRRRRR
RR
R--Ns00H0LkCCR8OsDNNF0HMFRVsHR#MCoDRk#FsROC8HC#oNMIsRC
RRRRRNRR0H0sLCk0RM#$_HLkDM0H_R8k:0R#soHM;R
RRRRRR0RN0LsHkR0C#_$MLDkH0_HM8FkRVWR7jb._s_F8#Rkl:MRC0$H0RRH#"NIC	
";RRRRRRRRRRRRRRRRRRRRRRRRRRRRS
SSCRM87.Wj_Fbs8k_#lR;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRS
SS
s
NO0EHCkO0ssCR0FDRVWR7jb._s_F8#RklH
#
-N-R0H0sLCk0RO8CDNNs0MHFRsVFRM#HoRDC#sFkO8CRCo#HMsINCRR
RRRRRNRR0H0sLCk0RM#$_HLkDM0H_R8k:0R#soHM;R
RRRRRR0RN0LsHkR0C#_$MLDkH0_HM8FkRV0RsDRR:NEsOHO0C0CksRRH#"NIC	
";
R--wRFs#oHMD#CRFOksCWR7,sRNO0EHCkO0s#CREDFk8CRLRl8klS$
Ns00H0LkC$R#MD_LN_O	LRFG:FRLFNDCMS;
Ns00H0LkC$R#MD_LN_O	LRFGFsVR0:DRRONsECH0Os0kC#RHRk0sC
;
LHCoM


CRM8s;0D
-
-============================================CHM00N$RMN8RsHOE00COkRsCVRFs8.Ij_OlN=============================D

HNLssQ$R ;  
Ck#R Q  03#8F_Do_HO4c4n3DND;#
kCCRHC#C30D8_FOoH_#kMHCoM8D3ND
;
CHM007$RW_j.lRNOHS#

MoCCOsH5S
SSIq_HE80Rh:Rq)azq=p:.R;
RRRRRRRRRARR_8IH0:ERRahqzp)q:
=4SRSRR;S2
bSSF5s0
SSSq:RSRRHM#_08DHFoOC_POs0F5Iq_HE80-84RF0IMF2Rj;S
SSSAR:MRHR8#0_oDFHPO_CFO0s_5AI0H8ER-48MFI0jFR2S;
SRSBSH:RM0R#8F_Do_HOP0COFqs5_8IH0+ERRIA_HE80-84RF0IMF2Rj;S
SSRaBSH:RM0R#8F_Do;HO
SSSvSqB:kRF00R#8F_Do_HOP0COFqs5_8IH0+ERRIA_HE80-84RF0IMF2Rj
SSS2-;
-0RN0LsHkR0C8DCON0sNHRFMVRFs#oHMD#CRFOksCCR8#MHoICNs
RRRRRRRR0N0skHL0#CR$LM_k0HDH8M_kRR:#H0sM
o;RRRRRRRRNs00H0LkC$R#Mk_LHHD0Mk_8RRFV7.Wj_OlNRC:RM00H$#RHRC"IN;	"
M
C8WR7jl._N
O;
ONsECH0Os0kC0RsDVRFRj7W.N_lO#RHS


-N-R0H0sLCk0RO8CDNNs0MHFRsVFRM#HoRDC#sFkO8CRCo#HMsINCRR
RRRRRNRR0H0sLCk0RM#$_HLkDM0H_R8k:0R#soHM;R
RRRRRR0RN0LsHkR0C#_$MLDkH0_HM8FkRV0RsDRR:NEsOHO0C0CksRRH#"NIC	
";
R--wRFs#oHMD#CRFOksCWR7,sRNO0EHCkO0s#CREDFk8CRLRl8klS$
Ns00H0LkC$R#MD_LN_O	LRFG:FRLFNDCMS;
Ns00H0LkC$R#MD_LN_O	LRFGFsVR0:DRRONsECH0Os0kC#RHRk0sC
;
LHCoM

SCRM8s;0D
-

-========================================C==M00H$MRN8sRNO0EHCkO0sVCRF8sRIH_8PC_sl=R======================R==
H
DLssN$ RQ 
 ;kR#CQ   38#0_oDFH4O_43ncN;DD
Ck#RCHCC03#8F_Do_HOkHM#o8MC3DND;#
kCCRHC#C30D8_FOoH_HNs0NE3D
D;
MSC0$H0R_7W8_HPsRClHS#
oCCMs5HO
SSSNH_I8R0E:1umQeaQ R:=US;
S_SLI0H8EuR:ma1QQ:e =;RU
SSS0lO_FR8C:aQh )t RR:=4SRS
SSS2S;
SsbF0S5
SRSNS:SSRRHM#_08DHFoOC_POs0F5IN_HE80-84RF0IMF2Rj;S
SSSLRSRS:H#MR0D8_FOoH_OPC05FsLH_I8-0E4FR8IFM0R;j2
SSS0SOSSH:RM0R#8F_Do;HO
SSSsNClHCM8sRS:FRk0#_08DHFoOC_POs0F5IL_HE80-84RF0IMF2Rj;S
SSFJk0MHC0RS:FRk0#_08DHFoOC_POs0F5IN_HE80-84RF0IMF2Rj;S
SSP8HH_8CLj$_SF:Rk#0R0D8_FOoH
SSS2-;
-0RN0LsHkR0C8DCON0sNHRFMVRFs#oHMD#CRFOksCCR8#MHoICNs
RRRRRRRR0N0skHL0#CR$LM_k0HDH8M_kRR:#H0sM
o;RRRRRRRRNs00H0LkC$R#Mk_LHHD0Mk_8RRFV78W_HsP_C:lRR0CMHR0$H"#RI	CN"
;
S8CMR_7W8_HPs;Cl
N

sHOE00COkRsCsR0DF7VRWH_8PC_sl#RHR-

-0RN0LsHkR0C8DCON0sNHRFMVRFs#oHMD#CRFOksCCR8#MHoICNsRR
RRRRRR0RN0LsHkR0C#_$MLDkH0_HM8:kRRs#0H;Mo
RRRRRRRR0N0skHL0#CR$LM_k0HDH8M_kVRFRDs0RN:RsHOE00COkRsCH"#RI	CN"
;
-w-RF#sRHDMoCFR#kCsOR,7WRONsECH0Os0kCER#F8kDRRLC8lkl$N
S0H0sLCk0RM#$_NLDOL	_F:GRRFLFDMCN;N
S0H0sLCk0RM#$_NLDOL	_FFGRV0RsDRR:NEsOHO0C0CksRRH#0Csk;S


LS
CMoH
M
C80RsD
;

=--=========================================0CMHR0$NRM8NEsOHO0C0CksRsVFRj7W.k_lD=0R========================
LDHs$NsR Q  k;
#QCR 3  #_08DHFoO4_4nNc3D
D;kR#CHCCC38#0_oDFHkO_Mo#HM3C8N;DD
Ck#RCHCC03#8F_Do_HON0sHED3ND
;

0CMHR0$7.Wj_Dlk0#RH
CSoMHCsO_5qI0H8EA,R_8IH0:ERR#bFHP0HC;R2
FSbs
05SRSqSRS:HSMR#_08DHFoOC_POs0F5IN_HE80-84RF0IMF2Rj;S
SASRS:MRHR0S#8F_Do_HOP0COFLs5_8IH04E-RI8FMR0Fj
2;SBSaR:SSRRHMS8#0_oDFH
O;S)SumB7zaRR:FRk0S8#0_oDFHPO_CFO0s_5NI0H8E_+LI0H8ER-48MFI0jFR2S
S2-;
-0RN0LsHkR0C8DCON0sNHRFMVRFs#oHMD#CRFOksCCR8#MHoICNs
RRRRRRRR0N0skHL0#CR$LM_k0HDH8M_kRR:#H0sM
o;RRRRRRRRNs00H0LkC$R#Mk_LHHD0Mk_8RRFV7.Wj_Dlk0RR:CHM00H$R#IR"C"N	;C

M78RW_j.l0kDR
;
NEsOHO0C0CksRDs0RRFV7.Wj_Dlk0#RHR-

-0RN0LsHkR0C8DCON0sNHRFMVRFs#oHMD#CRFOksCCR8#MHoICNsRR
RRRRRR0RN0LsHkR0C#_$MLDkH0_HM8:kRRs#0H;Mo
RRRRRRRR0N0skHL0#CR$LM_k0HDH8M_kVRFRDs0RN:RsHOE00COkRsCH"#RI	CN"
;
-w-RF#sRHDMoCFR#kCsOR,7WRONsECH0Os0kCER#F8kDRRLC8lkl$N
S0H0sLCk0RM#$_NLDOL	_F:GRRFLFDMCN;N
S0H0sLCk0RM#$_NLDOL	_FFGRV0RsDRR:NEsOHO0C0CksRRH#0Csk;L

CMoH
M
C80RsD
;
-=-=========================================CHM00N$RMN8RsHOE00COkRsCVRFs7.Wj_s#J0=R======================
==DsHLNRs$Q   ;#
kC RQ # 30D8_FOoH_n44cD3NDk;
#HCRC3CC#_08DHFoOM_k#MHoCN83D
D;kR#CHCCC38#0_oDFHNO_sEH03DND;C

M00H$WR7j#._JRs0Ho#
CsMCH
O5SISSHE80Su:Rma1QQRe :c=R;S
SS_aBlCF8RQ:Rhta  R)R:
=4S2SS;S
Sb0Fs5S
SS:qSRMRHR0S#8F_Do_HOP0COFIs5HE80-84RF0IMF2Rj;S
SSRaBRR:RHSMR#_08DHFoOS;
SmS)mRa:R0FkR0S#8F_Do_HOP0COF5s5I0H8E2+4/4.-RI8FMR0FjS2
S;S2
-
-R0N0skHL08CRCNODsHN0FVMRF#sRHDMoCFR#kCsOR#8CHIoMN
sCRRRRRRRRNs00H0LkC$R#Mk_LHHD0Mk_8R#:R0MsHoR;
RRRRRNRR0H0sLCk0RM#$_HLkDM0H_R8kF7VRW_j.#0JsRC:RM00H$#RHRC"IN;	"
M
C8WR7j#._J;s0
s
NO0EHCkO0ssCR0FDRVWR7j#._JRs0H
#
-N-R0H0sLCk0RO8CDNNs0MHFRsVFRM#HoRDC#sFkO8CRCo#HMsINCRR
RRRRRNRR0H0sLCk0RM#$_HLkDM0H_R8k:0R#soHM;R
RRRRRR0RN0LsHkR0C#_$MLDkH0_HM8FkRV0RsDRR:NEsOHO0C0CksRRH#"NIC	
";
R--wRFs#oHMD#CRFOksCWR7,sRNO0EHCkO0s#CREDFk8CRLRl8klS$
Ns00H0LkC$R#MD_LN_O	LRFG:FRLFNDCMS;
Ns00H0LkC$R#MD_LN_O	LRFGFsVR0:DRRONsECH0Os0kC#RHRk0sC
;
LHCoMC

Ms8R0
D;
=--=========================================0CMHR0$NRM8NEsOHO0C0CksRsVFR_7W1NJks=CR========================
LDHs$NsR Q  k;
#QCR 3  #_08DHFoO4_4nNc3D
D;kR#CQ   38#0_oDFHkO_Mo#HM3C8N;DD
C

M00H$WR7_k#JNRsCHo#
CsMCH
O5SHSI8R0E:qRhaqz)p4:=
2SS;b
SF5s0
NSSSRS:RRHMS8#0_oDFHPO_CFO0sH5I8-0E4FR8IFM0R;j2
0SSO:SSRMRHR0S#8F_Do;HOSS
S#NJks:CSRkRF0#RS0D8_FOoH_OPC05Fs5*.RR8IH0-E24FR8IFM0R
j2S;S2S-
-R0N0skHL08CRCNODsHN0FVMRF#sRHDMoCFR#kCsOR#8CHIoMN
sCRRRRRRRRNs00H0LkC$R#Mk_LHHD0Mk_8R#:R0MsHoR;
RRRRRNRR0H0sLCk0RM#$_HLkDM0H_R8kF7VRWJ_#kCNsRC:RM00H$#RHRC"IN;	"
M
C8WR7_k#JN;sC
s
NO0EHCkO0ssCR0FDRVWR7_k#JNRsCH-#
-0RN0LsHkR0C8DCON0sNHRFMVRFs#oHMD#CRFOksCCR8#MHoICNsRR
RRRRRR0RN0LsHkR0C#_$MLDkH0_HM8:kRRs#0H;Mo
RRRRRRRR0N0skHL0#CR$LM_k0HDH8M_kVRFRDs0RN:RsHOE00COkRsCH"#RI	CN"
;
-w-RF#sRHDMoCFR#kCsOR,7WRONsECH0Os0kCER#F8kDRRLC8lkl$N
S0H0sLCk0RM#$_NLDOL	_F:GRRFLFDMCN;N
S0H0sLCk0RM#$_NLDOL	_FFGRV0RsDRR:NEsOHO0C0CksRRH#0Csk;

RLHCoMC

Ms8R0RD;
-

-========================================C==M00H$MRN8sRNO0EHCkO0sVCRF7sRW_j.8HHP8=CR========================
H
DLssN$ RQ 
 ;kR#CQ   38#0_oDFH4O_43ncN;DD
Ck#RCHCC03#8F_Do_HOkHM#o8MC3DND;#
kCCRHC#C30D8_FOoH_HNs0NE3D
D;
0CMHR0$7.Wj_P8HHR8CH
#
oCCMs5HO
qSS_8IH0:ERR1umQeaQ =R:R
U;S_SAI0H8ERR:uQm1a QeRR:=US;
S_aBlCF8RQ:Rhta  :)R=
R4S;S2
FSbs
05SSSqSRS:HSMR#_08DHFoOC_POs0F5Iq_HE80-84RF0IMF2Rj;S
SASSS:MRHR0S#8F_Do_HOP0COFAs5_8IH04E-RI8FMR0Fj
2;SBSaS:SSRRHMS8#0_oDFH
O;SQS7e Q7__AYjRS:FRk0S8#0_oDFH
O;SzSTm aQh:aSR0FkR0S#8F_Do_HOP0COFqs5_8IH04E-RI8FMR0FjS2S
2SS;
SS-N-R0H0sLCk0RO8CDNNs0MHFRsVFRM#HoRDC#sFkO8CRCo#HMsINCR
RRRRRR0RN0LsHkR0C#_$MLDkH0_HM8:kRRs#0H;Mo
RRRRRRRR0N0skHL0#CR$LM_k0HDH8M_kVRFRj7W.H_8PCH8RC:RM00H$#RHRC"IN;	"
M
C8WR7j8._H8PHC
R;
ONsECH0Os0kC0RsDVRFRj7W.H_8PCH8RRH#
-
-R0N0skHL08CRCNODsHN0FVMRF#sRHDMoCFR#kCsOR#8CHIoMNRsC
RRRRRRRR0N0skHL0#CR$LM_k0HDH8M_kRR:#H0sM
o;RRRRRRRRNs00H0LkC$R#Mk_LHHD0Mk_8RRFVsR0D:sRNO0EHCkO0sHCR#IR"C"N	;-

-FRwsHR#MCoDRk#FsROC7RW,NEsOHO0C0CksRF#EkRD8L8CRk$ll
0SN0LsHkR0C#_$MLODN	F_LGRR:LDFFC;NM
0SN0LsHkR0C#_$MLODN	F_LGVRFRDs0RN:RsHOE00COkRsCH0#Rs;kC
L

CMoH
M
C80RsD
;

=--============================================CHM00N$RMN8RsHOE00COkRsCVRFs7PW_Cls_F=8R========================
LDHs$NsR Q  k;
#QCR 3  #_08DHFoO4_4nNc3D
D;kR#CHCCC38#0_oDFHkO_Mo#HM3C8N;DD
Ck#RCHCC03#8F_Do_HON0sHED3ND
;
CHM007$RWC_PsF_l8#RH
C
oMHCsOS5
SIq_HE80Ru:Rma1QQRe :c=R;S
SAH_I8R0E:mRu1QQae: R=;R.
aSSBF_l8:CRRaQh )t R=R:RS4
S
2;SsbF0S5
SSqS:HRRM#RS0D8_FOoH_OPC05FsqH_I8-0E4FR8IFM0R;j2
ASSSRS:RRHMS8#0_oDFHPO_CFO0s_5AI0H8ER-48MFI0jFR2S;
SSaBSR:RHSMR#_08DHFoOS;
S7vmz1pzSR:RFRk0S8#0_oDFHPO_CFO0s_5AI0H8ER-48MFI0jFR2S
S2-;
-0RN0LsHkR0C8DCON0sNHRFMVRFs#oHMD#CRFOksCCR8#MHoICNs
RRRRRRRR0N0skHL0#CR$LM_k0HDH8M_kRR:#H0sM
o;RRRRRRRRNs00H0LkC$R#Mk_LHHD0Mk_8RRFV7PW_Cls_F:8RR0CMHR0$H"#RI	CN"
;
 RM87PW_Cls_F;8R
s
NO0EHCkO0ssCR0FDRVWR7_sPC_8lFRRH#
-
-R0N0skHL08CRCNODsHN0FVMRF#sRHDMoCFR#kCsOR#8CHIoMNRsC
RRRRRRRR0N0skHL0#CR$LM_k0HDH8M_kRR:#H0sM
o;RRRRRRRRNs00H0LkC$R#Mk_LHHD0Mk_8RRFVsR0D:sRNO0EHCkO0sHCR#IR"C"N	;-

-FRwsHR#MCoDRk#FsROC7RW,NEsOHO0C0CksRF#EkRD8L8CRk$ll
0SN0LsHkR0C#_$MLODN	F_LGRR:LDFFC;NM
0SN0LsHkR0C#_$MLODN	F_LGVRFRDs0RN:RsHOE00COkRsCH0#Rs;kC
L

CMoH
M
C80RsD
;
-=-==========================================C==M00H$MRN8sRNO0EHCkO0sVCRF7sRW_j.sRCl=========================H
DLssN$ RQ 
 ;kR#CQ   38#0_oDFH4O_43ncN;DD
Ck#RCHCC03#8F_Do_HOkHM#o8MC3DND;#
kCCRHC#C30D8_FOoH_HNs0NE3D
D;
0CMHR0$7.Wj_lsCR
H#
MoCCOsH5S
SqH_I8R0E:mRu1QQae: R=;R.
ASS_8IH0:ERR1umQeaQ =R:R
.;SBSa_8lFCRR:Q hatR )RR:=4S
S2S;
b0Fs5S
SqSSS:HRRM#RS0D8_FOoH_OPC05FsqH_I8-0E4FR8IFM0R;j2
ASSS:SSRMRHR0S#8F_Do_HOP0COFAs5_8IH04E-RI8FMR0Fj
2;SBSaS:SSRMRHR0S#8F_Do;HO
)SS Qvqh)7 SR:RFRk0S8#0_oDFHPO_CFO0s_5AI0H8ER-48MFI0jFR2S
S2S;R
R--Ns00H0LkCCR8OsDNNF0HMFRVsHR#MCoDRk#FsROC8HC#oNMIsRC
RRRRRNRR0H0sLCk0RM#$_HLkDM0H_R8k:0R#soHM;R
RRRRRR0RN0LsHkR0C#_$MLDkH0_HM8FkRVWR7js._C:lRR0CMHR0$H"#RI	CN"
;
CRM87.Wj_lsCR
;
NEsOHO0C0CksRDs0RRFV7.Wj_lsCRRH#
-
-R0N0skHL08CRCNODsHN0FVMRF#sRHDMoCFR#kCsOR#8CHIoMNRsC
RRRRRRRR0N0skHL0#CR$LM_k0HDH8M_kRR:#H0sM
o;RRRRRRRRNs00H0LkC$R#Mk_LHHD0Mk_8RRFVsR0D:sRNO0EHCkO0sHCR#IR"C"N	;-

-FRwsHR#MCoDRk#FsROC7RW,NEsOHO0C0CksRF#EkRD8L8CRk$ll
0SN0LsHkR0C#_$MLODN	F_LGRR:LDFFC;NM
0SN0LsHkR0C#_$MLODN	F_LGVRFRDs0RN:RsHOE00COkRsCH0#Rs;kC


SS

SLHCoMC

Ms8R0
D;
=--============================================CHM00N$RMN8RsHOE00COkRsCVRFs7eW_]l7_F=8R========================
LDHs$NsR Q  k;
#QCR 3  #_08DHFoO4_4nNc3D
D;kR#CHCCC38#0_oDFHkO_Mo#HM3C8N;DD
Ck#RCHCC03#8F_Do_HON0sHED3ND
;
CHM007$RWE_P8F_l8#RH
MoCCOsH5S
SqH_I8R0E:mRu1QQae: R=;Rc
ASS_8IH0:ERR1umQeaQ =R:R
d;SBSa_8lFCRR:Q hatR )RR:=4S
S2S;
b0Fs5S
SqSRRSR:RHSMR#_08DHFoOC_POs0F5Iq_HE80-84RF0IMF2Rj;S
SASRRSR:RHSMR#_08DHFoOC_POs0F5IA_HE80-84RF0IMF2Rj;S
SaSBRSR:RHSMR#_08DHFoOS;
S7vmz1pzRR:RFRk0S8#0_oDFHPO_CFO0s_5AI0H8ER-48MFI0jFR2S
S2
;S-N-R0H0sLCk0RO8CDNNs0MHFRsVFRM#HoRDC#sFkO8CRCo#HMsINCR
RRRRRR0RN0LsHkR0C#_$MLDkH0_HM8:kRRs#0H;Mo
RRRRRRRR0N0skHL0#CR$LM_k0HDH8M_kVRFR_7WP_E8lRF8:MRC0$H0RRH#"NIC	
";
8CMR_7WP_E8lRF8;N

sHOE00COkRsCsR0DF7VRWE_P8F_l8#RH
-
-R0N0skHL08CRCNODsHN0FVMRF#sRHDMoCFR#kCsOR#8CHIoMNRsC
RRRRRRRR0N0skHL0#CR$LM_k0HDH8M_kRR:#H0sM
o;RRRRRRRRNs00H0LkC$R#Mk_LHHD0Mk_8RRFVsR0D:sRNO0EHCkO0sHCR#IR"C"N	;-

-FRwsHR#MCoDRk#FsROC7RW,NEsOHO0C0CksRF#EkRD8L8CRk$ll
0SN0LsHkR0C#_$MLODN	F_LGRR:LDFFC;NM
0SN0LsHkR0C#_$MLODN	F_LGVRFRDs0RN:RsHOE00COkRsCH0#Rs;kC
SR

oLCH
M
CRM8s;0D
