library verilog;
use verilog.vl_types.all;
entity MRRST_N_TREE is
    port(
        A               : in     vl_logic;
        Z               : out    vl_logic
    );
end MRRST_N_TREE;
