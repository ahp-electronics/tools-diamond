library verilog;
use verilog.vl_types.all;
entity PCNTR_delc1x2v1s is
    port(
        A               : in     vl_logic;
        Z               : out    vl_logic
    );
end PCNTR_delc1x2v1s;
