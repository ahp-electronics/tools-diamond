library verilog;
use verilog.vl_types.all;
entity ebr_hse_top is
    port(
        addr_1          : in     vl_logic;
        addr_0          : in     vl_logic;
        cib_addra_12    : in     vl_logic;
        cib_addra_11    : in     vl_logic;
        cib_addra_10    : in     vl_logic;
        cib_addra_9     : in     vl_logic;
        cib_addra_8     : in     vl_logic;
        cib_addra_7     : in     vl_logic;
        cib_addra_6     : in     vl_logic;
        cib_addra_5     : in     vl_logic;
        cib_addra_4     : in     vl_logic;
        cib_addra_3     : in     vl_logic;
        cib_addra_2     : in     vl_logic;
        cib_addra_1     : in     vl_logic;
        cib_addra_0     : in     vl_logic;
        cib_addrb_12    : in     vl_logic;
        cib_addrb_11    : in     vl_logic;
        cib_addrb_10    : in     vl_logic;
        cib_addrb_9     : in     vl_logic;
        cib_addrb_8     : in     vl_logic;
        cib_addrb_7     : in     vl_logic;
        cib_addrb_6     : in     vl_logic;
        cib_addrb_5     : in     vl_logic;
        cib_addrb_4     : in     vl_logic;
        cib_addrb_3     : in     vl_logic;
        cib_addrb_2     : in     vl_logic;
        cib_addrb_1     : in     vl_logic;
        cib_addrb_0     : in     vl_logic;
        cib_cea         : in     vl_logic;
        cib_ceb         : in     vl_logic;
        cib_clka        : in     vl_logic;
        cib_clkb        : in     vl_logic;
        cib_csa_2       : in     vl_logic;
        cib_csa_1       : in     vl_logic;
        cib_csa_0       : in     vl_logic;
        cib_csb_2       : in     vl_logic;
        cib_csb_1       : in     vl_logic;
        cib_csb_0       : in     vl_logic;
        cib_dataa_8     : in     vl_logic;
        cib_dataa_7     : in     vl_logic;
        cib_dataa_6     : in     vl_logic;
        cib_dataa_5     : in     vl_logic;
        cib_dataa_4     : in     vl_logic;
        cib_dataa_3     : in     vl_logic;
        cib_dataa_2     : in     vl_logic;
        cib_dataa_1     : in     vl_logic;
        cib_dataa_0     : in     vl_logic;
        cib_datab_8     : in     vl_logic;
        cib_datab_7     : in     vl_logic;
        cib_datab_6     : in     vl_logic;
        cib_datab_5     : in     vl_logic;
        cib_datab_4     : in     vl_logic;
        cib_datab_3     : in     vl_logic;
        cib_datab_2     : in     vl_logic;
        cib_datab_1     : in     vl_logic;
        cib_datab_0     : in     vl_logic;
        cib_oprcea      : in     vl_logic;
        cib_oprceb      : in     vl_logic;
        cib_rsta        : in     vl_logic;
        cib_rstb        : in     vl_logic;
        cib_wea         : in     vl_logic;
        cib_web         : in     vl_logic;
        es_o_35         : in     vl_logic;
        es_o_34         : in     vl_logic;
        es_o_33         : in     vl_logic;
        es_o_32         : in     vl_logic;
        es_o_31         : in     vl_logic;
        es_o_30         : in     vl_logic;
        es_o_29         : in     vl_logic;
        es_o_28         : in     vl_logic;
        es_o_27         : in     vl_logic;
        es_o_26         : in     vl_logic;
        es_o_25         : in     vl_logic;
        es_o_24         : in     vl_logic;
        es_o_23         : in     vl_logic;
        es_o_22         : in     vl_logic;
        es_o_21         : in     vl_logic;
        es_o_20         : in     vl_logic;
        es_o_19         : in     vl_logic;
        es_o_18         : in     vl_logic;
        es_o_17         : in     vl_logic;
        es_o_16         : in     vl_logic;
        es_o_15         : in     vl_logic;
        es_o_14         : in     vl_logic;
        es_o_13         : in     vl_logic;
        es_o_12         : in     vl_logic;
        es_o_11         : in     vl_logic;
        es_o_10         : in     vl_logic;
        es_o_9          : in     vl_logic;
        es_o_8          : in     vl_logic;
        es_o_7          : in     vl_logic;
        es_o_6          : in     vl_logic;
        es_o_5          : in     vl_logic;
        es_o_4          : in     vl_logic;
        es_o_3          : in     vl_logic;
        es_o_2          : in     vl_logic;
        es_o_1          : in     vl_logic;
        es_o_0          : in     vl_logic;
        from_prev_ebr_8 : in     vl_logic;
        from_prev_ebr_7 : in     vl_logic;
        from_prev_ebr_6 : in     vl_logic;
        from_prev_ebr_5 : in     vl_logic;
        from_prev_ebr_4 : in     vl_logic;
        from_prev_ebr_3 : in     vl_logic;
        from_prev_ebr_2 : in     vl_logic;
        from_prev_ebr_1 : in     vl_logic;
        from_prev_ebr_0 : in     vl_logic;
        from_prev_sel   : in     vl_logic;
        gsrn            : in     vl_logic;
        por_n           : in     vl_logic;
        trim_mem_2      : in     vl_logic;
        trim_mem_1      : in     vl_logic;
        trim_mem_0      : in     vl_logic;
        vccm            : in     vl_logic;
        aempty_flag     : out    vl_logic;
        afull_flag      : out    vl_logic;
        doa_8           : out    vl_logic;
        doa_7           : out    vl_logic;
        doa_6           : out    vl_logic;
        doa_5           : out    vl_logic;
        doa_4           : out    vl_logic;
        doa_3           : out    vl_logic;
        doa_2           : out    vl_logic;
        doa_1           : out    vl_logic;
        doa_0           : out    vl_logic;
        dob_8           : out    vl_logic;
        dob_7           : out    vl_logic;
        dob_6           : out    vl_logic;
        dob_5           : out    vl_logic;
        dob_4           : out    vl_logic;
        dob_3           : out    vl_logic;
        dob_2           : out    vl_logic;
        dob_1           : out    vl_logic;
        dob_0           : out    vl_logic;
        empty_flag      : out    vl_logic;
        full_flag       : out    vl_logic;
        mc1_out_39      : out    vl_logic;
        mc1_out_38      : out    vl_logic;
        mc1_out_37      : out    vl_logic;
        mc1_out_36      : out    vl_logic;
        mc1_out_35      : out    vl_logic;
        mc1_out_34      : out    vl_logic;
        mc1_out_33      : out    vl_logic;
        mc1_out_32      : out    vl_logic;
        mc1_out_31      : out    vl_logic;
        mc1_out_30      : out    vl_logic;
        mc1_out_29      : out    vl_logic;
        mc1_out_28      : out    vl_logic;
        mc1_out_27      : out    vl_logic;
        mc1_out_26      : out    vl_logic;
        mc1_out_25      : out    vl_logic;
        mc1_out_24      : out    vl_logic;
        mc1_out_23      : out    vl_logic;
        mc1_out_22      : out    vl_logic;
        mc1_out_21      : out    vl_logic;
        mc1_out_20      : out    vl_logic;
        mc1_out_19      : out    vl_logic;
        mc1_out_18      : out    vl_logic;
        mc1_out_17      : out    vl_logic;
        mc1_out_16      : out    vl_logic;
        mc1_out_15      : out    vl_logic;
        mc1_out_14      : out    vl_logic;
        mc1_out_13      : out    vl_logic;
        mc1_out_12      : out    vl_logic;
        mc1_out_11      : out    vl_logic;
        mc1_out_10      : out    vl_logic;
        mc1_out_9       : out    vl_logic;
        mc1_out_8       : out    vl_logic;
        mc1_out_7       : out    vl_logic;
        mc1_out_6       : out    vl_logic;
        mc1_out_5       : out    vl_logic;
        mc1_out_4       : out    vl_logic;
        mc1_out_3       : out    vl_logic;
        mc1_out_2       : out    vl_logic;
        mc1_out_1       : out    vl_logic;
        mc1_out_0       : out    vl_logic;
        to_next_ebr_8   : out    vl_logic;
        to_next_ebr_7   : out    vl_logic;
        to_next_ebr_6   : out    vl_logic;
        to_next_ebr_5   : out    vl_logic;
        to_next_ebr_4   : out    vl_logic;
        to_next_ebr_3   : out    vl_logic;
        to_next_ebr_2   : out    vl_logic;
        to_next_ebr_1   : out    vl_logic;
        to_next_ebr_0   : out    vl_logic;
        to_next_sel     : out    vl_logic;
        data_143        : inout  vl_logic;
        data_142        : inout  vl_logic;
        data_141        : inout  vl_logic;
        data_140        : inout  vl_logic;
        data_139        : inout  vl_logic;
        data_138        : inout  vl_logic;
        data_137        : inout  vl_logic;
        data_136        : inout  vl_logic;
        data_135        : inout  vl_logic;
        data_134        : inout  vl_logic;
        data_133        : inout  vl_logic;
        data_132        : inout  vl_logic;
        data_131        : inout  vl_logic;
        data_130        : inout  vl_logic;
        data_129        : inout  vl_logic;
        data_128        : inout  vl_logic;
        data_127        : inout  vl_logic;
        data_126        : inout  vl_logic;
        data_125        : inout  vl_logic;
        data_124        : inout  vl_logic;
        data_123        : inout  vl_logic;
        data_122        : inout  vl_logic;
        data_121        : inout  vl_logic;
        data_120        : inout  vl_logic;
        data_119        : inout  vl_logic;
        data_118        : inout  vl_logic;
        data_117        : inout  vl_logic;
        data_116        : inout  vl_logic;
        data_115        : inout  vl_logic;
        data_114        : inout  vl_logic;
        data_113        : inout  vl_logic;
        data_112        : inout  vl_logic;
        data_111        : inout  vl_logic;
        data_110        : inout  vl_logic;
        data_109        : inout  vl_logic;
        data_108        : inout  vl_logic;
        data_107        : inout  vl_logic;
        data_106        : inout  vl_logic;
        data_105        : inout  vl_logic;
        data_104        : inout  vl_logic;
        data_103        : inout  vl_logic;
        data_102        : inout  vl_logic;
        data_101        : inout  vl_logic;
        data_100        : inout  vl_logic;
        data_99         : inout  vl_logic;
        data_98         : inout  vl_logic;
        data_97         : inout  vl_logic;
        data_96         : inout  vl_logic;
        data_95         : inout  vl_logic;
        data_94         : inout  vl_logic;
        data_93         : inout  vl_logic;
        data_92         : inout  vl_logic;
        data_91         : inout  vl_logic;
        data_90         : inout  vl_logic;
        data_89         : inout  vl_logic;
        data_88         : inout  vl_logic;
        data_87         : inout  vl_logic;
        data_86         : inout  vl_logic;
        data_85         : inout  vl_logic;
        data_84         : inout  vl_logic;
        data_83         : inout  vl_logic;
        data_82         : inout  vl_logic;
        data_81         : inout  vl_logic;
        data_80         : inout  vl_logic;
        data_79         : inout  vl_logic;
        data_78         : inout  vl_logic;
        data_77         : inout  vl_logic;
        data_76         : inout  vl_logic;
        data_75         : inout  vl_logic;
        data_74         : inout  vl_logic;
        data_73         : inout  vl_logic;
        data_72         : inout  vl_logic;
        data_71         : inout  vl_logic;
        data_70         : inout  vl_logic;
        data_69         : inout  vl_logic;
        data_68         : inout  vl_logic;
        data_67         : inout  vl_logic;
        data_66         : inout  vl_logic;
        data_65         : inout  vl_logic;
        data_64         : inout  vl_logic;
        data_63         : inout  vl_logic;
        data_62         : inout  vl_logic;
        data_61         : inout  vl_logic;
        data_60         : inout  vl_logic;
        data_59         : inout  vl_logic;
        data_58         : inout  vl_logic;
        data_57         : inout  vl_logic;
        data_56         : inout  vl_logic;
        data_55         : inout  vl_logic;
        data_54         : inout  vl_logic;
        data_53         : inout  vl_logic;
        data_52         : inout  vl_logic;
        data_51         : inout  vl_logic;
        data_50         : inout  vl_logic;
        data_49         : inout  vl_logic;
        data_48         : inout  vl_logic;
        data_47         : inout  vl_logic;
        data_46         : inout  vl_logic;
        data_45         : inout  vl_logic;
        data_44         : inout  vl_logic;
        data_43         : inout  vl_logic;
        data_42         : inout  vl_logic;
        data_41         : inout  vl_logic;
        data_40         : inout  vl_logic;
        data_39         : inout  vl_logic;
        data_38         : inout  vl_logic;
        data_37         : inout  vl_logic;
        data_36         : inout  vl_logic;
        data_35         : inout  vl_logic;
        data_34         : inout  vl_logic;
        data_33         : inout  vl_logic;
        data_32         : inout  vl_logic;
        data_31         : inout  vl_logic;
        data_30         : inout  vl_logic;
        data_29         : inout  vl_logic;
        data_28         : inout  vl_logic;
        data_27         : inout  vl_logic;
        data_26         : inout  vl_logic;
        data_25         : inout  vl_logic;
        data_24         : inout  vl_logic;
        data_23         : inout  vl_logic;
        data_22         : inout  vl_logic;
        data_21         : inout  vl_logic;
        data_20         : inout  vl_logic;
        data_19         : inout  vl_logic;
        data_18         : inout  vl_logic;
        data_17         : inout  vl_logic;
        data_16         : inout  vl_logic;
        data_15         : inout  vl_logic;
        data_14         : inout  vl_logic;
        data_13         : inout  vl_logic;
        data_12         : inout  vl_logic;
        data_11         : inout  vl_logic;
        data_10         : inout  vl_logic;
        data_9          : inout  vl_logic;
        data_8          : inout  vl_logic;
        data_7          : inout  vl_logic;
        data_6          : inout  vl_logic;
        data_5          : inout  vl_logic;
        data_4          : inout  vl_logic;
        data_3          : inout  vl_logic;
        data_2          : inout  vl_logic;
        data_1          : inout  vl_logic;
        data_0          : inout  vl_logic;
        datan_143       : inout  vl_logic;
        datan_142       : inout  vl_logic;
        datan_141       : inout  vl_logic;
        datan_140       : inout  vl_logic;
        datan_139       : inout  vl_logic;
        datan_138       : inout  vl_logic;
        datan_137       : inout  vl_logic;
        datan_136       : inout  vl_logic;
        datan_135       : inout  vl_logic;
        datan_134       : inout  vl_logic;
        datan_133       : inout  vl_logic;
        datan_132       : inout  vl_logic;
        datan_131       : inout  vl_logic;
        datan_130       : inout  vl_logic;
        datan_129       : inout  vl_logic;
        datan_128       : inout  vl_logic;
        datan_127       : inout  vl_logic;
        datan_126       : inout  vl_logic;
        datan_125       : inout  vl_logic;
        datan_124       : inout  vl_logic;
        datan_123       : inout  vl_logic;
        datan_122       : inout  vl_logic;
        datan_121       : inout  vl_logic;
        datan_120       : inout  vl_logic;
        datan_119       : inout  vl_logic;
        datan_118       : inout  vl_logic;
        datan_117       : inout  vl_logic;
        datan_116       : inout  vl_logic;
        datan_115       : inout  vl_logic;
        datan_114       : inout  vl_logic;
        datan_113       : inout  vl_logic;
        datan_112       : inout  vl_logic;
        datan_111       : inout  vl_logic;
        datan_110       : inout  vl_logic;
        datan_109       : inout  vl_logic;
        datan_108       : inout  vl_logic;
        datan_107       : inout  vl_logic;
        datan_106       : inout  vl_logic;
        datan_105       : inout  vl_logic;
        datan_104       : inout  vl_logic;
        datan_103       : inout  vl_logic;
        datan_102       : inout  vl_logic;
        datan_101       : inout  vl_logic;
        datan_100       : inout  vl_logic;
        datan_99        : inout  vl_logic;
        datan_98        : inout  vl_logic;
        datan_97        : inout  vl_logic;
        datan_96        : inout  vl_logic;
        datan_95        : inout  vl_logic;
        datan_94        : inout  vl_logic;
        datan_93        : inout  vl_logic;
        datan_92        : inout  vl_logic;
        datan_91        : inout  vl_logic;
        datan_90        : inout  vl_logic;
        datan_89        : inout  vl_logic;
        datan_88        : inout  vl_logic;
        datan_87        : inout  vl_logic;
        datan_86        : inout  vl_logic;
        datan_85        : inout  vl_logic;
        datan_84        : inout  vl_logic;
        datan_83        : inout  vl_logic;
        datan_82        : inout  vl_logic;
        datan_81        : inout  vl_logic;
        datan_80        : inout  vl_logic;
        datan_79        : inout  vl_logic;
        datan_78        : inout  vl_logic;
        datan_77        : inout  vl_logic;
        datan_76        : inout  vl_logic;
        datan_75        : inout  vl_logic;
        datan_74        : inout  vl_logic;
        datan_73        : inout  vl_logic;
        datan_72        : inout  vl_logic;
        datan_71        : inout  vl_logic;
        datan_70        : inout  vl_logic;
        datan_69        : inout  vl_logic;
        datan_68        : inout  vl_logic;
        datan_67        : inout  vl_logic;
        datan_66        : inout  vl_logic;
        datan_65        : inout  vl_logic;
        datan_64        : inout  vl_logic;
        datan_63        : inout  vl_logic;
        datan_62        : inout  vl_logic;
        datan_61        : inout  vl_logic;
        datan_60        : inout  vl_logic;
        datan_59        : inout  vl_logic;
        datan_58        : inout  vl_logic;
        datan_57        : inout  vl_logic;
        datan_56        : inout  vl_logic;
        datan_55        : inout  vl_logic;
        datan_54        : inout  vl_logic;
        datan_53        : inout  vl_logic;
        datan_52        : inout  vl_logic;
        datan_51        : inout  vl_logic;
        datan_50        : inout  vl_logic;
        datan_49        : inout  vl_logic;
        datan_48        : inout  vl_logic;
        datan_47        : inout  vl_logic;
        datan_46        : inout  vl_logic;
        datan_45        : inout  vl_logic;
        datan_44        : inout  vl_logic;
        datan_43        : inout  vl_logic;
        datan_42        : inout  vl_logic;
        datan_41        : inout  vl_logic;
        datan_40        : inout  vl_logic;
        datan_39        : inout  vl_logic;
        datan_38        : inout  vl_logic;
        datan_37        : inout  vl_logic;
        datan_36        : inout  vl_logic;
        datan_35        : inout  vl_logic;
        datan_34        : inout  vl_logic;
        datan_33        : inout  vl_logic;
        datan_32        : inout  vl_logic;
        datan_31        : inout  vl_logic;
        datan_30        : inout  vl_logic;
        datan_29        : inout  vl_logic;
        datan_28        : inout  vl_logic;
        datan_27        : inout  vl_logic;
        datan_26        : inout  vl_logic;
        datan_25        : inout  vl_logic;
        datan_24        : inout  vl_logic;
        datan_23        : inout  vl_logic;
        datan_22        : inout  vl_logic;
        datan_21        : inout  vl_logic;
        datan_20        : inout  vl_logic;
        datan_19        : inout  vl_logic;
        datan_18        : inout  vl_logic;
        datan_17        : inout  vl_logic;
        datan_16        : inout  vl_logic;
        datan_15        : inout  vl_logic;
        datan_14        : inout  vl_logic;
        datan_13        : inout  vl_logic;
        datan_12        : inout  vl_logic;
        datan_11        : inout  vl_logic;
        datan_10        : inout  vl_logic;
        datan_9         : inout  vl_logic;
        datan_8         : inout  vl_logic;
        datan_7         : inout  vl_logic;
        datan_6         : inout  vl_logic;
        datan_5         : inout  vl_logic;
        datan_4         : inout  vl_logic;
        datan_3         : inout  vl_logic;
        datan_2         : inout  vl_logic;
        datan_1         : inout  vl_logic;
        datan_0         : inout  vl_logic
    );
end ebr_hse_top;
