library verilog;
use verilog.vl_types.all;
entity ebr_hse_fusebox is
    port(
        vccm            : inout  vl_logic;
        vssm            : inout  vl_logic;
        addr            : in     vl_logic_vector(1 downto 0);
        data            : inout  vl_logic_vector(143 downto 0);
        datan           : inout  vl_logic_vector(143 downto 0);
        es_mode         : in     vl_logic;
        f_unused        : out    vl_logic_vector(39 downto 0);
        f_wta           : out    vl_logic;
        f_wtb           : out    vl_logic;
        f_rbwa          : out    vl_logic;
        f_rbwb          : out    vl_logic;
        f_mfg_mem       : out    vl_logic_vector(10 downto 0);
        f_doublewidea   : out    vl_logic;
        f_w_ctrl_a      : out    vl_logic_vector(2 downto 0);
        f_doublewideb   : out    vl_logic;
        f_w_ctrl_b      : out    vl_logic_vector(2 downto 0);
        f_wid           : out    vl_logic_vector(8 downto 0);
        f_rid           : out    vl_logic_vector(8 downto 0);
        f_wen           : out    vl_logic_vector(1 downto 0);
        f_ren           : out    vl_logic;
        f_oregsela      : out    vl_logic;
        f_oregselb      : out    vl_logic;
        async_fuse      : out    vl_logic;
        f_grdis         : out    vl_logic;
        f_ebr_enable    : out    vl_logic;
        f_pcsa          : out    vl_logic_vector(2 downto 0);
        f_pcsb          : out    vl_logic_vector(2 downto 0);
        f_prsta         : out    vl_logic;
        f_prstb         : out    vl_logic;
        f_pw_ra         : out    vl_logic;
        f_pw_rb         : out    vl_logic;
        f_n_edge        : out    vl_logic;
        f_mfg_spc       : out    vl_logic_vector(4 downto 0);
        f_spc           : out    vl_logic;
        f_addra         : out    vl_logic_vector(1 downto 0);
        f_addra_p       : out    vl_logic_vector(1 downto 0);
        f_addrb_0       : out    vl_logic;
        f_addrb_p_0     : out    vl_logic;
        f_mfg_clka      : out    vl_logic_vector(1 downto 0);
        f_mfg_clkb      : out    vl_logic_vector(1 downto 0);
        f_rst_sync_dis  : out    vl_logic;
        f_fifo_en       : out    vl_logic;
        f_pf            : out    vl_logic_vector(13 downto 0);
        f_pfm1          : out    vl_logic_vector(13 downto 0);
        f_paf           : out    vl_logic_vector(13 downto 0);
        f_pafm1         : out    vl_logic_vector(13 downto 0);
        f_1shot         : out    vl_logic;
        f_min_delay     : out    vl_logic;
        f_max_delay     : out    vl_logic;
        f_e             : out    vl_logic_vector(4 downto 0);
        f_ep1           : out    vl_logic_vector(5 downto 0);
        f_pae           : out    vl_logic_vector(13 downto 0);
        f_paep1         : out    vl_logic_vector(13 downto 0);
        fifo_rdw        : out    vl_logic_vector(2 downto 0);
        fifo_wdw        : out    vl_logic_vector(2 downto 0)
    );
end ebr_hse_fusebox;
