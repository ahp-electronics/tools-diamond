library verilog;
use verilog.vl_types.all;
entity UM_DEL is
    port(
        A               : in     vl_logic;
        Y               : out    vl_logic
    );
end UM_DEL;
