library verilog;
use verilog.vl_types.all;
entity cdr_alu is
    generic(
        STATE_INI       : integer := 0;
        STATE_ADD       : integer := 1;
        STATE_RUN       : integer := 3;
        STATE_FDN       : integer := 2
    );
    port(
        L0              : out    vl_logic_vector(3 downto 0);
        L1              : out    vl_logic_vector(3 downto 0);
        L2              : out    vl_logic_vector(3 downto 0);
        L3              : out    vl_logic_vector(3 downto 0);
        L4              : out    vl_logic_vector(3 downto 0);
        L5              : out    vl_logic_vector(3 downto 0);
        L6              : out    vl_logic_vector(3 downto 0);
        L7              : out    vl_logic_vector(3 downto 0);
        L8              : out    vl_logic_vector(3 downto 0);
        L9              : out    vl_logic_vector(3 downto 0);
        L10             : out    vl_logic_vector(3 downto 0);
        L11             : out    vl_logic_vector(3 downto 0);
        L12             : out    vl_logic_vector(3 downto 0);
        L13             : out    vl_logic_vector(3 downto 0);
        L14             : out    vl_logic_vector(3 downto 0);
        L15             : out    vl_logic_vector(3 downto 0);
        L16             : out    vl_logic_vector(3 downto 0);
        L17             : out    vl_logic_vector(3 downto 0);
        M0              : out    vl_logic_vector(3 downto 0);
        M1              : out    vl_logic_vector(3 downto 0);
        M2              : out    vl_logic_vector(3 downto 0);
        M3              : out    vl_logic_vector(3 downto 0);
        M4              : out    vl_logic_vector(3 downto 0);
        M5              : out    vl_logic_vector(3 downto 0);
        M6              : out    vl_logic_vector(3 downto 0);
        M7              : out    vl_logic_vector(3 downto 0);
        M8              : out    vl_logic_vector(3 downto 0);
        M9              : out    vl_logic_vector(3 downto 0);
        M10             : out    vl_logic_vector(3 downto 0);
        M11             : out    vl_logic_vector(3 downto 0);
        M12             : out    vl_logic_vector(3 downto 0);
        M13             : out    vl_logic_vector(3 downto 0);
        M14             : out    vl_logic_vector(3 downto 0);
        M15             : out    vl_logic_vector(3 downto 0);
        M16             : out    vl_logic_vector(3 downto 0);
        M17             : out    vl_logic_vector(3 downto 0);
        START_LOCK      : out    vl_logic;
        ACLK            : in     vl_logic;
        SEL_WIDTH       : in     vl_logic;
        CR0             : in     vl_logic;
        CR1             : in     vl_logic;
        CR2             : in     vl_logic;
        CR3             : in     vl_logic;
        CR4             : in     vl_logic;
        CR5             : in     vl_logic;
        CR6             : in     vl_logic;
        CR7             : in     vl_logic;
        CR8             : in     vl_logic;
        CR9             : in     vl_logic;
        CR10            : in     vl_logic;
        CR11            : in     vl_logic;
        CR12            : in     vl_logic;
        CR13            : in     vl_logic;
        CR14            : in     vl_logic;
        CR15            : in     vl_logic;
        CR16            : in     vl_logic;
        CR17            : in     vl_logic;
        RST_N           : in     vl_logic;
        LOCK            : in     vl_logic;
        UP_DN           : in     vl_logic;
        HOLD_ALU        : in     vl_logic;
        MC1_BW          : in     vl_logic_vector(1 downto 0)
    );
end cdr_alu;
