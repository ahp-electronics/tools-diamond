--
@ER--B$FbsEHo0OR52gR4g-cRRj.jd$R1MHbDO$H0ROQM
R--fN]C8:CsR#//$DMbH0OH$N/lb..jjDjdNl0/NCbbsN#/0D0/HoL/CFM_sdONON/sl__sIE3P8Ry4f-
-
-

--
-

---7-Rk-NDb0FsRv)qR0IHECR#bNCs0qCR7 7)1V1RFssRCRN8NRM8I0sHC-
-RsaNoRC0:kRpO0CMRm-R)RBqd-B
-H
DLssN$CRHC
C;kR#CHCCC38#0_oDFH4O_43ncN;DD
Ck#RCHCC03#8F_Do_HO#MHoCN83D
D;kR#CHCCC38#0_oDFHNO_sEH03DND;H
DLssN$sRFO;Nd
Ck#ROFsNFd3sOONF3lbN;DD
0CMHR0$)_qv)R_WHR#
RoRRCsMCH5OR
RRRRRRRRlVNH:D$Rs#0HRMo:"=RMCFM"R;
RRRRRIRRHE80RH:RMo0CC:sR=;R(RR
RRRRRR8RN8HsI8R0E:MRH0CCos=R:RR(;RRRRR-RR-HRLoMRCFEkoRsVFRb8C0RE
RRRRR8RRCEb0RH:RMo0CC:sR=4RR.
U;RRRRRRRR80Fk_osCRL:RFCFDN:MR=NRVD;#CRRRRRR--ERN#Fbk0ks0RCRo
RRRRR8RRHsM_C:oRRFLFDMCNRR:=V#NDCR;RRRRR-E-RN8#RNR0NHkMb0CRsoR
RRRRRRNRs8_8ssRCo:FRLFNDCM=R:RDVN#RC;R-RR-NRE8CRsNN8R8C8s#s#RCRo
RRRRRIRRNs88_osCRL:RFCFDN:MR=NRVDR#CRRRR-E-RNI8RsCH0R8N8s#C#RosC
RRRRRRRR
2;RRRRb0FsRR5
RRRRR7RRmRzaRF:Rk#0R0D8_FOoH_OPC05FsI0H8ER-48MFI0jFR2R;
RRRRR)RRq)77RH:RM#RR0D8_FOoH_OPC05FsNs88I0H8ER-48MFI0jFR2R;
RRRRR7RRQRhRRH:RM#RR0D8_FOoH_OPC05FsI0H8ER-48MFI0jFR2R;
RRRRRWRRq)77RH:RM#RR0D8_FOoH_OPC05FsNs88I0H8ER-48MFI0jFR2R;
RRRRRWRR RRRRH:RM#RR0D8_FOoH;RRRRRRR-I-RsCH0RNCMLRDCVRFss
NlRRRRRRRRBRpiRRR:HRMR#_08DHFoOR;RRRRRRR--OODF	FRVsNRslN,R8,8sRM8H
RRRRRRRRpmBi:RRRRHMR8#0_oDFHRORRRRRR-R-R0FbRFODOV	RF8sRF
k0RRRRRRRR2C;
MC8RM00H$qR)v__)W
;
---
-HRwsR#0HDlbCMlC0HN0FlMRkR#0LOCRNCDD8sRNO
Ej-N-
sHOE00COkRsCNEsOjVRFRv)q_W)_R
H#O#FM00NMRlMk_DOCD8#_CRCb:MRH0CCos=R:R855CEb0R4-R2./d2R;RRRRRR-RR-RRyFsVRFRI#F7VRB. dXOcRC#DDRCMC8
C8O#FM00NMRlMk_DOCDI#_HR8C:MRH0CCos=R:RI55HE80R4-R22/c;RRRRRRRR-RR-RRyFOVRFlDkMF#RVBR7 Xd.cCRODRD#M8CCC08
$RbCF_k0L_k#0C$bRRH#NNss$MR5kOl_C#DD_C8CbFR8IFM0RRj,5lMk_DOCDI#_H*8Ccd2+RI8FMR0FjF2RV0R#8F_Do;HO
o#HMRNDF_k0LRk#:kRF0k_L#$_0bRC;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-.-R7sRNsRN$F8VRFRk05bHMk00RFsR0H0-#N#0C2H
#oDMNR0Fk_RCMR:RRR8#0_oDFHPO_CFO0sk5MlC_OD_D#8bCCRI8FMR0FjR2;RR--CLMNDRC#VRFs0-sH#00NC##
HNoMDbRICCj_MRRR:0R#8F_Do_HOP0COFMs5kOl_C#DD_C8CbFR8IFM0R;j2R-R-RHIs0CCRMDNLCV#RFCsRNROEsRFIF)VRqOvRC#DD
o#HMRNDI4bC_RCMRRR:#_08DHFoOC_POs0F5lMk_DOCD8#_CRCb8MFI0jFR2R;R-I-RsCH0RNCML#DCRsVFROCNEFRsIVRFRv)qRDOCD##
HNoMDMRH_osCRRRR:0R#8F_Do_HOP0COFIs5HE80+8dRF0IMF2Rj;RRRRRRRR-R-RCk#8FR0RosCHC#0sQR7h#R
HNoMD RW_t) 4RRR:0R#8F_Do;HO
o#HMRNDHsM_CRo4RRR:#_08DHFoOC_POs0F58IH0dE+RI8FMR0FjR2;R
RR#MHoNFDRks0_CRoRR#:R0D8_FOoH_OPC05FsI0H8ER+d8MFI0jFR2R;RRRRRR-RR-#RkC08RFCRso0H#C7sRm
za#MHoNsDRNs8_CRoRR#:R0D8_FOoH_OPC05FsNs88I0H8ER-48MFI0jFR2R;RR-RR-#RkC08RFCRso0H#C)sRq)77
o#HMRNDI_N8sRCoRRR:#_08DHFoOC_POs0F58N8s8IH04E-RI8FMR0FjR2;RRRR-k-R#RC80sFRC#oH0RCsW7q7)H
#oDMNRIDF_8sN8:sRR8#0_oDFHPO_CFO0sR5c8MFI0jFR2R;RRRRRRRRRRRRRRR--s8N8sHRL0H#RM0bkRR0F)RqvODCD#6R5R0LH#CRsJskHC
82#MHoNDDRFII_Ns88R#:R0D8_FOoH_OPC05FscFR8IFM0R;j2RRRRRRRRRRRRR-RR-NRI8R8sL#H0RbHMk00RFqR)vCRODRD#5L6RHR0#skCJH8sC2$
0b0CRlNb_8_8s0C$bRRH#NNss$MR5kOl_C#DD_C8CbFR8IFM0RRj2F#VR0D8_FOoH_OPC0RFs58gRF0IMF2Rj;H
#oDMNRb0l_8N8s:RRRb0l_8N8s$_0b
C;
oLCH
M
RRRR-Q-RV8RN8HsI8R0E<RR6NH##o'MRj0'RFMRkk8#CR0LH#R
RR4RzRRR:H5VRNs88I0H8ERR=4o2RCsMCN
0CRRRRRRRRD_FIs8N8s=R<Rj"jjRj"&NRs8C_so25j;R
RRRRRRFRDIN_I8R8s<"=Rjjjj"RR&I_N8s5Coj
2;RRRRCRM8oCCMsCN0R;z4
RRRRRz.RH:RVNR58I8sHE80R.=R2CRoMNCs0RC
RRRRRDRRFsI_Ns88RR<="jjj"RR&s_N8s5Co4FR8IFM0R;j2
RRRRRRRRIDF_8IN8<sR=jR"jRj"&NRI8C_soR548MFI0jFR2R;
RCRRMo8RCsMCNR0Cz
.;RRRRzRdR:VRHR85N8HsI8R0E=2RdRMoCC0sNCR
RRRRRRFRDIN_s8R8s<"=RjRj"&NRs8C_soR5.8MFI0jFR2R;
RRRRRDRRFII_Ns88RR<=""jjRI&RNs8_C.o5RI8FMR0Fj
2;RRRRCRM8oCCMsCN0R;zd
RRRRRzcRH:RVNR58I8sHE80Rc=R2CRoMNCs0RC
RRRRRDRRFsI_Ns88RR<='Rj'&NRs8C_soR5d8MFI0jFR2R;
RRRRRDRRFII_Ns88RR<='Rj'&NRI8C_soR5d8MFI0jFR2R;
RCRRMo8RCsMCNR0Cz
c;RRRRzR6R:VRHR85N8HsI8R0E>2RcRMoCC0sNCR
RRRRRRFRDIN_s8R8s<s=RNs8_Cco5RI8FMR0Fj
2;RRRRRRRRD_FII8N8s=R<R8IN_osC58cRF0IMF2Rj;R
RRMRC8CRoMNCs0zCR6
;
RRRR-Q-RV8R5HsM_CRo2sHCo#s0CRh7QRHk#MBoRpRi
RzRRn:RRRRHV5M8H_osC2CRoMNCs0RC
RRRRRbRRsCFO#5#RB,piRh7Q2CRLo
HMRRRRRRRRRRRRH5VRBRpi=4R''MRN8pRBiP'CC2M0RC0EMR
RRRRRRRRRRRRRRMRH_osCRR<=5j"jjRj"&QR7h
2;RRRRRRRRRRRRCRM8H
V;RRRRRRRRCRM8bOsFC;##
RRRR8CMRMoCC0sNCnRz;R
RR(RzRRR:H5VRMRF08_HMs2CoRMoCC0sNCR
RRRRRRRRRRMRH_osCRR<=5j"jjRj"&QR7h
2;RRRRCRM8oCCMsCN0R;z(
R
RR-R-RRQV58sN8ss_CRo2sHCo#s0CR7)q7k)R#oHMRiBp
RRRRjz4RRR:H5VRs8N8sC_soo2RCsMCN
0CRRRRRRRRbOsFCR##5pmBi),Rq)772CRLo
HMRRRRRRRRRRRRH5VRmiBpR'=R4N'RMm8RB'piCMPC002RE
CMRRRRRRRRRRRRRRRRs_N8sRCo<)=Rq)7758N8s8IH04E-RI8FMR0Fj
2;RRRRRRRRRRRRCRM8H
V;RRRRRRRRCRM8bOsFC;##
RRRR8CMRMoCC0sNC4RzjR;
RzRR4:4RRRHV50MFR8sN8ss_CRo2oCCMsCN0
RRRRRRRRRRRR8sN_osCRR<=)7q7)85N8HsI8-0E4FR8IFM0R;j2
RRRR8CMRMoCC0sNC4Rz4R;
RRRRR
RRRRRR-Q-RVIR5Ns88_osC2CRso0H#CWsRq)77RHk#MBoRpRi
RzRR4R.R:VRHRN5I8_8ss2CoRMoCC0sNCR
RRRRRRsRbF#OC#BR5pRi,W7q7)L2RCMoH
RRRRRRRRRRRRRHV5iBpR'=R4N'RMB8RpCi'P0CM2ER0CRM
RRRRRRRRRRRRRIRRNs8_C<oR=qRW757)Ns88I0H8ER-48MFI0jFR2R;
RRRRRRRRRCRRMH8RVR;
RRRRRCRRMb8RsCFO#
#;RRRRCRM8oCCMsCN0R.z4;R
RR4RzdRR:H5VRMRF0I8N8sC_soo2RCsMCN
0CRRRRRRRRRRRRI_N8sRCo<W=Rq)77;R
RRMRC8CRoMNCs0zCR4
d;
RRRRR--tCCMsCN0RC0ERv)qRDOCDN#RM#8RCODC0FRDo
HORRRRzR4c:FRVsRRHHMMRkOl_C#DD_C8CbFR8IFM0RojRCsMCN
0CRRRR-A-Rk8HDR0FkbRk0CLMND#CRCODC0FRDo
HORRRRRRRR-Q-RVNR58I8sHE80R4>R6O2RN0M'RCk#R1NRpRQBODCD
RRRRRRRR4m nRR:H5VRNs88I0H8ERR>4R62oCCMsCN0
RRRRRRRRRRRRRRRR0Fk_5CMH<2R=4R''ERIC5MRs_N8s5CoNs88I0H8ER-48MFI06FR2RR=HC2RDR#C';j'
RRRRRRRR8CMRMoCC0sNC Rm4
n;RRRRRRRR-Q-RVNR58I8sHE80R6>R2hRq7NR58I8sHE80RR<=4R62kR#NNpR1QOBRC
DDRRRRRRRRm6 4RH:RVNR58I8sHE80R4=R6o2RCsMCN
0CRRRRRRRRRRRRRRRR0_lbNs8855H2gFR8IFM0RRj2<h=RmOa5F_MP#_08DHFoOC_POs0F5RH,42j2R)XmR8sN_osC58N8s8IH04E-RI8FMR0F6
2;RRRRRRRRRRRRRRRR17qh_R46:qR1hj74RsbF0NRlbqR5RR=>0_lbNs8855H2jR2,A>R=Rb0l_8N8s25H5,42R=BR>lR0b8_N8Hs5225.,RR7=0>RlNb_858sHd252R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR =0>RlNb_858sHc252w,RRR=>0_lbNs8855H26R2,t>R=Rb0l_8N8s25H5,n2R=]R>lR0b8_N8Hs5225(,RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRQ=0>RlNb_858sHU252K,RRR=>0_lbNs8855H2gR2,Z>R=R0Fk_5CMH;22
RRRRRRRR8CMRMoCC0sNC Rm4
6;RRRRRRRRmc 4RH:RVNR58I8sHE80R4=Rco2RCsMCN
0CRRRRRRRRRRRRRRRR0_lbNs8855H2UFR8IFM0RRj2<h=RmOa5F_MP#_08DHFoOC_POs0F5RH,gR22XRm)s_N8s5CoNs88I0H8ER-48MFI06FR2R;
RRRRRRRRRRRRR1RRq_h74:cRRh1q7R4jb0FsRblNRR5q=0>RlNb_858sHj252A,RRR=>0_lbNs8855H24R2,B>R=Rb0l_8N8s25H5,.2R=7R>lR0b8_N8Hs5225d,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR= R>lR0b8_N8Hs5225c,RRw=0>RlNb_858sH6252t,RRR=>0_lbNs8855H2nR2,]>R=Rb0l_8N8s25H5,(2RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR=QR>lR0b8_N8Hs5225U,RRK='>R4R',Z>R=R0Fk_5CMH;22
RRRRRRRR8CMRMoCC0sNC Rm4
c;RRRRRRRRmd 4RH:RVNR58I8sHE80R4=Rdo2RCsMCN
0CRRRRRRRRRRRRRRRR0_lbNs8855H2(FR8IFM0RRj2<h=RmOa5F_MP#_08DHFoOC_POs0F5RH,UR22XRm)s_N8s5CoNs88I0H8ER-48MFI06FR2R;
RRRRRRRRRRRRR1RRq_h74:dRRh1q7RURb0FsRblNRR5q=0>RlNb_858sHj252A,RRR=>0_lbNs8855H24R2,B>R=Rb0l_8N8s25H5,.2R=7R>lR0b8_N8Hs5225d,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR= R>lR0b8_N8Hs5225c,RRw=0>RlNb_858sH6252t,RRR=>0_lbNs8855H2nR2,]>R=Rb0l_8N8s25H5,(2RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR=ZR>kRF0M_C52H2;R
RRRRRRMRC8CRoMNCs0mCR ;4d
RRRRRRRR4m .RR:H5VRNs88I0H8ERR=4R.2oCCMsCN0
RRRRRRRRRRRRRRRRb0l_8N8s25H58nRF0IMF2RjRR<=h5maOPFM_8#0_oDFHPO_CFO0s,5HR2(2R)XmR8sN_osC58N8s8IH04E-RI8FMR0F6
2;RRRRRRRRRRRRRRRR17qh_R4.:qR1hR7URsbF0NRlbqR5RR=>0_lbNs8855H2jR2,A>R=Rb0l_8N8s25H5,42R=BR>lR0b8_N8Hs5225.,RR7=0>RlNb_858sHd252R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR =0>RlNb_858sHc252w,RRR=>0_lbNs8855H26R2,t>R=Rb0l_8N8s25H5,n2R=]R>4R''
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRZRRRR=>F_k0CHM52
2;RRRRRRRRCRM8oCCMsCN0R4m .R;
RRRRRmRR R44:VRHR85N8HsI8R0E=4R42CRoMNCs0RC
RRRRRRRRRRRRR0RRlNb_858sH625RI8FMR0Fj<2R=mRhaF5OM#P_0D8_FOoH_OPC05FsHn,R2X2Rms)RNs8_CNo58I8sHE80-84RF0IMF2R6;R
RRRRRRRRRRRRRRqR1h47_4RR:17qhnbRRFRs0lRNb5=qR>lR0b8_N8Hs5225j,RRA=0>RlNb_858sH4252B,RRR=>0_lbNs8855H2.R2,7>R=Rb0l_8N8s25H5,d2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR >R=Rb0l_8N8s25H5,c2R=wR>lR0b8_N8Hs52256,RRZ=F>RkC0_M25H2R;
RRRRRCRRMo8RCsMCNR0Cm4 4;R
RRRRRR Rm4:jRRRHV58N8s8IH0=ERR24jRMoCC0sNCR
RRRRRRRRRRRRRRlR0b8_N8Hs52R5c8MFI0jFR2=R<Rahm5MOFP0_#8F_Do_HOP0COFHs5,2R62mRX)NRs8C_so85N8HsI8-0E4FR8IFM0R;62
RRRRRRRRRRRRRRRRh1q7j_4R1:Rqnh7RFRbsl0RN5bRq>R=Rb0l_8N8s25H5,j2R=AR>lR0b8_N8Hs52254,RRB=0>RlNb_858sH.2527,RRR=>0_lbNs8855H2d
2,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR RRRR=>0_lbNs8855H2cR2,w>R=R''4,RRZ=F>RkC0_M25H2R;
RRRRRCRRMo8RCsMCNR0Cmj 4;R
RRRRRR Rmg:RRRRHV58N8s8IH0=ERRRg2oCCMsCN0
RRRRRRRRRRRRRRRRb0l_8N8s25H58dRF0IMF2RjRR<=h5maOPFM_8#0_oDFHPO_CFO0s,5HR2c2R)XmR8sN_osC58N8s8IH04E-RI8FMR0F6
2;RRRRRRRRRRRRRRRR17qh_:gRRh1q7RcRRsbF0NRlbqR5RR=>0_lbNs8855H2jR2,A>R=Rb0l_8N8s25H5,42R=BR>lR0b8_N8Hs5225.,RR7=0>RlNb_858sHd252R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRZ=F>RkC0_M25H2R;
RRRRRCRRMo8RCsMCNR0Cm; g
RRRRRRRRUm RRR:H5VRNs88I0H8ERR=Uo2RCsMCN
0CRRRRRRRRRRRRRRRR0_lbNs8855H2.FR8IFM0RRj2<h=RmOa5F_MP#_08DHFoOC_POs0F5RH,dR22XRm)s_N8s5CoNs88I0H8ER-48MFI06FR2R;
RRRRRRRRRRRRR1RRq_h7URR:17qhcRRRb0FsRblNRR5q=0>RlNb_858sHj252A,RRR=>0_lbNs8855H24R2,B>R=Rb0l_8N8s25H5,.2R=7R>4R''R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRZ=F>RkC0_M25H2R;
RRRRRCRRMo8RCsMCNR0Cm; U
RRRRRRRR(m RRR:H5VRNs88I0H8ERR=(o2RCsMCN
0CRRRRRRRRRRRRRRRR0_lbNs8855H24FR8IFM0RRj2<h=RmOa5F_MP#_08DHFoOC_POs0F5RH,.R22XRm)s_N8s5CoNs88I0H8ER-48MFI06FR2R;
RRRRRRRRRRRRR1RRq_h7(RR:17qh.RRRb0FsRblNRR5q=0>RlNb_858sHj252A,RRR=>0_lbNs8855H24R2,Z>R=R0Fk_5CMH;22
RRRRRRRR8CMRMoCC0sNC Rm(R;
RRRRRmRR RnR:VRHR85N8HsI8R0E=2RnRMoCC0sNCR
RRRRRRRRRRRRRRkRF0M_C5RH2<'=R4I'RERCM58sN_osC5R62=FROM#P_0D8_FOoH_OPC05FsH2,452j2R#CDCjR''R;
RRRRRCRRMo8RCsMCNR0Cm; n
RRRRR--Q5VRNs88I0H8E=R<RR62MFFRkk0b0MRCNCLDRD#CCRO0DHFoOCRMC88C
RRRRRRRR6m RH:RVNR58I8sHE80RR<=6o2RCsMCN
0CRRRRRRRRRRRRRRRRF_k0CHM52=R<R''4;R
RRRRRRMRC8CRoMNCs0mCR 
6;
RRRRR--Q5VRNs88I0H8ERR>gk2R#WCRuR j08FRC8OFC8RN8#sC#HRL0n#RRs0EFEkoRNgRMW8RuR 408FRC8OFCHRL04#Rj
R+RRRRRRRRWj 4RH:RVNR58I8sHE80Rg>R2CRoMNCs0RC
RRRRRRRRRRRRRIRRb_CjCHM52=R<R''4RCIEMIR5Ns8_CUo5RI8FMR0F6=2RRMOFP0_#8F_Do_HOP0COFHs5,2.j58dRF0IMF2Rj2DRC#'CRj
';RRRRRRRRRRRRRRRRI4bC_5CMH<2R=4R''ERIC5MRI_N8s5CoNs88I0H8ER-48MFI0gFR2RR=OPFM_8#0_oDFHPO_CFO0s,5H.5j2Ns88I0H8ER-n8MFI0cFR2C2RDR#C';j'
RRRRRRRRRRRR8CMRMoCC0sNC RW4
j;RRRR-Q-RVNR58I8sHE80RU=RRRFsgk2R#WCRuR j08FRC8OFC8RN8#sC#HRL0n#RRs0EFEkoRRg
RRRRRWRR RgR:VRHRN558I8sHE80RU=R2)RmR85N8HsI8R0E=2Rg2CRoMNCs0RC
RRRRRRRRRRRRRIRRb_CjCHM52=R<R''4RCIEMIR5Ns8_CNo58I8sHE80-84RF0IMF2R6RH=R2DRC#'CRj
';RRRRRRRRRRRRRRRRI4bC_5CMH<2R=4R''R;
RRRRRRRRRCRRMo8RCsMCNR0CW; g
RRRRR--Q5VRNs88I0H8ERR=(k2R#WCRuR j08FRC8OFCER0C0RnE8RN8#sC#HRL0RR&W4u RR0F8FCO80CRE(CR0NER8C8s#L#RHR0
RRRRRWRR R(R:VRHR85N8HsI8R0E=2R(RMoCC0sNCR
RRRRRRRRRRRRRRbRICCj_M25HRR<='R4'IMECRN5I8C_so256RO=RF_MP#_08DHFoOC_POs0F5.H,225j2DRC#'CRj
';RRRRRRRRRRRRRRRRI4bC_5CMH<2R=4R''ERIC5MRI_N8s5Con=2RRMOFP0_#8F_Do_HOP0COFHs5,5.24R22CCD#R''j;R
RRRRRRMRC8CRoMNCs0WCR 
(;RRRR-Q-RVNR58I8sHE80Rn=R2#RkCuRW 0jRFCR8OCF8RC0EREn0R8N8s#C#R0LH
RRRRRRRRnW RRR:H5VRNs88I0H8ERR=no2RCsMCN
0CRRRRRRRRRRRRRRRRIjbC_5CMH<2R=4R''ERIC5MRI_N8s5Co6=2RRMOFP0_#8F_Do_HOP0COFHs5,542jR22CCD#R''j;R
RRRRRRRRRRRRRRbRICC4_M25HRR<=';4'
RRRRRRRR8CMRMoCC0sNC RWnR;
R-RR-VRQR85N8HsI8R0E<6=R2FRMRHIs0CCRMDNLCCR#D0CORoDFHMORCCC88R
RRRRRR RW6:RRRRHV58N8s8IH0<ER=2R6RMoCC0sNCR
RRRRRRRRRRRRRRbRICCj_M25HRR<=';4'
RRRRRRRRRRRRRRRRCIb4M_C5RH2<'=R4
';RRRRRRRRCRM8oCCMsCN0R6W ;R

RCRRMo8RCsMCNR0Cz;4c
R
RRsRbF#OC#BR5pRi,72QhRoLCHRM
RRRRRVRHRp5BiRR='R4'NRM8B'piCMPC002RE
CMRRRRRRRRRHRRMC_so<4R=MRH_osC;R
RRRRRRRRRR_W )4 tRR<=W
 ;RRRRRCRRMH8RVR;
RCRRMb8RsCFO#
#;
RRRR6z.RH:RVMR5F80RF_k0s2CoRMoCC0sNCR
RRRRRR4Rz(R4:bOsFCR##5_W )4 t,qR)7,7)R7Wq7R),HsM_C,o4R0Fk_osC2R
RRRRRRCRLo
HMRRRRRRRRRRRRH5VR5_W )4 tR'=R4R'2NRM857)q7=)RR7Wq72)2RC0EMR
RRRRRRRRRRRRRRmR7z<aR=MRH_osC4H5I8-0E4FR8IFM0R;j2
RRRRRRRRRRRR#CDCR
RRRRRRRRRRRRRRmR7z<aR=kRF0C_soH5I8-0E4FR8IFM0R;j2
RRRRRRRRRRRR8CMR;HV
RRRRRRRR8CMRFbsO#C#R(z44R;
RCRRMo8RCsMCNR0Cz;.6
R
RRdRzj:RRRRHV5k8F0C_soo2RCsMCN
0CRRRRRRRRbOsFCR##5pmBiF,Rks0_CRo2LHCoMR
RRRRRRRRRRVRHRB5mp=iRR''4R8NMRpmBiP'CC2M0RC0EMR
RRRRRRRRRRRRRRmR7z<aR=kRF0C_soH5I8-0E4FR8IFM0R;j2
RRRRRRRRRRRR8CMR;HV
RRRRRRRR8CMRFbsO#C#;R
RRMRC8CRoMNCs0zCRd
j;
RRRRR--tsMCNR0C0REC)RqvODCD#HRI00ERs#H-0CN0#R
RR4Rz6RR:VRFsHMRHRlMk_DOCD8#_CRCb8MFI0jFRRMoCC0sNCR
RRRRRR4Rz(RR:VRFs[MRHRlMk_DOCDI#_HR8C8MFI0jFRRMoCC0sNCR
RRRRRRRRRR)RzqRv:7dB .RXc
RRRRRRRRRRRRRRRRsbF0NRlb7R5Q=jR>MRH_osC5*5[c,22R47QRR=>HsM_C5o5[2*c+,42R.7QRR=>HsM_C5o5[2*c+,.2Rd7QRR=>HsM_C5o5[2*c+,d2
RRRRRRRRRRRRRRRRRRRRRRRRWRRqR7j=D>RFII_Ns885,j2R7Wq4>R=RIDF_8IN84s52W,RqR7.=D>RFII_Ns885,.2R7Wqd>R=RIDF_8IN8ds52W,RqR7c=D>RFII_Ns885,c2
RRRRRRRRRRRRRRRRRRRRRRRR)RRqR7j=D>RFsI_Ns885,j2R7)q4>R=RIDF_8sN84s52),RqR7.=D>RFsI_Ns885,.2R7)qd>R=RIDF_8sN8ds52),RqR7c=D>RFsI_Ns885,c2
R--RRRRRRRRRRRRRRRRRRRRRRRRR W)h>R=R,W R Wuj>R=RCIbjM_C5,H2R Wu4>R=RCIb4M_C5,H2RRBi=h>RmBa5p,i2RR
RRRRRRRRRRRRRRRRRRRRRRRRRWh) RR=>WR ,Wju RR=>IjbC_5CMHR2,W4u RR=>I4bC_5CMHR2,B=iR>pRBi
,RRRRRRRRRRRRRRRRRRRRRRRRRRmR7j>R=R0Fk_#Lk55H,[2*c27,Rm=4R>kRF0k_L#,5H5c[*22+4,mR7.>R=R0Fk_#Lk55H,[2*c+,.2Rd7mRR=>F_k0L5k#H[,5*+c2d;22
RRRRRRRRRRRRRRRR0Fk_osC5*5[cR22<F=RkL0_kH#5,*5[cR22IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*5[c42+2=R<R0Fk_#Lk55H,[2*c+R42IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*5[c.2+2=R<R0Fk_#Lk55H,[2*c+R.2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*5[cd2+2=R<R0Fk_#Lk55H,[2*c+Rd2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRR8CMRMoCC0sNC4Rz(R;
RCRRMo8RCsMCNR0Cz;46
-
-R.RzURR:H5VR80Fk_osC2CRoMNCs0-C
-RRRRRRRRnz4RV:RFHsRRRHMM_klODCD#C_8C8bRF0IMFRRjoCCMsCN0
R--RRRRRzRR4:URRsVFRH[RMkRMlC_OD_D#ICH8RI8FMR0FjCRoMNCs0-C
-RRRRRRRRRRRRqz)v7:RB. dX
cR-R-RRRRRRRRRRRRRRFRbsl0RN5bR7RQj=H>RMC_so[55*2c2,QR74>R=R_HMs5Co5c[*22+4,QR7.>R=R_HMs5Co5c[*22+.,QR7d>R=R_HMs5Co5c[*22+d,-
-RRRRRRRRRRRRRRRRRRRRRRRRRqRW7=jR>FRDIN_I858sjR2,W4q7RR=>D_FII8N8s254,qRW7=.R>FRDIN_I858s.R2,Wdq7RR=>D_FII8N8s25d,qRW7=cR>FRDIN_I858sc
2,-R-RRRRRRRRRRRRRRRRRRRRRRRRR)jq7RR=>D_FIs8N8s25j,qR)7=4R>FRDIN_s858s4R2,).q7RR=>D_FIs8N8s25.,qR)7=dR>FRDIN_s858sdR2,)cq7RR=>D_FIs8N8s25c,-
-RRRRRRRRRRRRRRRRRRRRRRRRR)RW =hR> RW,uRW =jR>bRICCj_M25H,uRW =4R>bRICC4_M25H,iRBRR=>h5maB2pi,-R
-RRRRRRRRRRRRRRRRRRRRRRRRTRR7Rmj=F>RkL0_kH#5,*5[c,22RmT74>R=R0Fk_#Lk55H,[2*c+,42RmT7.>R=R0Fk_#Lk55H,[2*c+,.2RmT7d>R=R0Fk_#Lk55H,[2*c+2d2;-
-
R--RRRRRRRRRRRRR0Fk_osC5*5[cR22<F=RkL0_kH#5,*5[cR22IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
R--RRRRRRRRRRRRRFRRks0_C5o5[2*c+R42<F=RkL0_kH#5,*5[c42+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''-;
-RRRRRRRRRRRRRRRR0Fk_osC5*5[c.2+2=R<R0Fk_#Lk55H,[2*c+R.2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
R--RRRRRRRRRRRRRFRRks0_C5o5[2*c+Rd2<F=RkL0_kH#5,*5[cd2+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''-;
-RRRRRRRRRRRR8CMRMoCC0sNC4RzU-;
-RRRRRRRCRM8oCCMsCN0Rnz4;-
-RRRRCRM8oCCMsCN0RUz.;-

-RRRRkRRURR:H5VR80Fk_osC2CRoMNCs0-C
-RRRR7RRmRza<F=Rks0_CIo5HE80-84RF0IMF2Rj;-
-RMRC8CRoMNCs0kCRUR;
RRRRR
RRCRM8NEsOHO0C0CksRONsE
j;
