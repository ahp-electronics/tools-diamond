library verilog;
use verilog.vl_types.all;
entity cfg_qual is
    port(
        jump_exec       : out    vl_logic;
        chip_select_exec: out    vl_logic;
        flow_through_exec: out    vl_logic;
        bypass_exec     : out    vl_logic;
        isc_data_shift_iqual: out    vl_logic;
        lsc_prog_incr_rti_iqual: out    vl_logic;
        lsc_prog_incr_enc_iqual: out    vl_logic;
        lsc_prog_incr_cmp_iqual: out    vl_logic;
        lsc_prog_incr_cne_iqual: out    vl_logic;
        isc_data_shift_cqual: out    vl_logic;
        lsc_prog_incr_rti_cqual: out    vl_logic;
        lsc_prog_incr_enc_cqual: out    vl_logic;
        lsc_prog_incr_cmp_cqual: out    vl_logic;
        lsc_prog_incr_cne_cqual: out    vl_logic;
        verify_id_qual  : out    vl_logic;
        read_temp_qual  : out    vl_logic;
        lsc_device_ctrl_qual: out    vl_logic;
        prog_dryrun_addr_qual: out    vl_logic;
        lsc_shift_password_qual: out    vl_logic;
        lsc_bitstream_burst_qual: out    vl_logic;
        sf_address_shift_qual: out    vl_logic;
        lsc_prog_ctrl0_qual: out    vl_logic;
        lsc_read_ctrl0_qual: out    vl_logic;
        lsc_prog_ctrl1_qual: out    vl_logic;
        lsc_read_ctrl1_qual: out    vl_logic;
        lsc_reset_crc_qual: out    vl_logic;
        lsc_read_crc_qual: out    vl_logic;
        lsc_write_comp_dic_qual: out    vl_logic;
        lsc_read_comp_dic_qual: out    vl_logic;
        sed_init_addr_qual: out    vl_logic;
        sed_write_addr_qual: out    vl_logic;
        sed_read_incr_qual: out    vl_logic;
        sed_prog_sed_crc_qual: out    vl_logic;
        sed_prog_ctrl0_qual: out    vl_logic;
        sed_prog_ctrl1_qual: out    vl_logic;
        sed_write_comp_dic_qual: out    vl_logic;
        sf_prog_ucode_qual: out    vl_logic;
        sf_program_qual : out    vl_logic;
        sf_read_qual    : out    vl_logic;
        sf_erase_qual   : out    vl_logic;
        sf_prog_done_qual: out    vl_logic;
        sf_erase_done_qual: out    vl_logic;
        sf_prog_sec_qual: out    vl_logic;
        sf_init_addr_qual: out    vl_logic;
        sf_write_addr_qual: out    vl_logic;
        sf_prog_incr_rti_qual: out    vl_logic;
        sf_prog_incr_enc_qual: out    vl_logic;
        sf_prog_incr_cmp_qual: out    vl_logic;
        sf_prog_incr_cne_qual: out    vl_logic;
        sf_vfy_incr_rti_qual: out    vl_logic;
        sf_prog_sed_crc_qual: out    vl_logic;
        sf_read_sed_crc_qual: out    vl_logic;
        sf_write_bus_addr_qual: out    vl_logic;
        sf_pcs_write_qual: out    vl_logic;
        sf_pcs_read_qual: out    vl_logic;
        sf_ebr_write_qual: out    vl_logic;
        sf_ebr_read_qual: out    vl_logic;
        sf_prog_sec_eqv : out    vl_logic;
        fl_erase_qual_pre: out    vl_logic;
        fl_prog_done_qual: out    vl_logic;
        fl_prog_sec_qual: out    vl_logic;
        fl_prog_secplus_qual: out    vl_logic;
        fl_prog_ucode_qual: out    vl_logic;
        fl_prog_authmode_qual: out    vl_logic;
        fl_prog_aesfea_qual: out    vl_logic;
        fl_init_addr_qual: out    vl_logic;
        fl_write_addr_qual: out    vl_logic;
        fl_prog_incr_nv_qual: out    vl_logic;
        fl_read_incr_nv_qual: out    vl_logic;
        fl_prog_password_qual: out    vl_logic;
        fl_prog_cipher_key0_qual: out    vl_logic;
        fl_prog_cipher_key1_qual: out    vl_logic;
        fl_prog_feature_qual: out    vl_logic;
        fl_prog_feabits_qual: out    vl_logic;
        fl_init_addr_ufm_qual: out    vl_logic;
        fl_prog_tag_qual: out    vl_logic;
        fl_erase_tag_qual: out    vl_logic;
        fl_read_tag_qual: out    vl_logic;
        fl_prog_pes_qual: out    vl_logic;
        fl_prog_mes_qual: out    vl_logic;
        fl_prog_hes_qual: out    vl_logic;
        fl_prog_trim0_qual: out    vl_logic;
        fl_prog_trim1_qual: out    vl_logic;
        fl_read_hes_qual: out    vl_logic;
        fl_prog_csec_qual: out    vl_logic;
        fl_prog_usec_qual: out    vl_logic;
        fl_prog_uds_qual: out    vl_logic;
        fl_mtest_qual   : out    vl_logic;
        mfg_margin_en   : out    vl_logic;
        mfg_flash_en    : out    vl_logic;
        dryrun_prog_ucode_qual: out    vl_logic;
        isc_prog_done_qual: out    vl_logic;
        isc_prog_sec_qual: out    vl_logic;
        isc_prog_secplus_qual: out    vl_logic;
        isc_prog_ucode_qual: out    vl_logic;
        lsc_prog_authdone0_qual: out    vl_logic;
        lsc_prog_authdone1_qual: out    vl_logic;
        lsc_prog_authmode_qual: out    vl_logic;
        lsc_prog_aesfea_qual: out    vl_logic;
        lsc_prog_password_qual: out    vl_logic;
        lsc_prog_cipher_key0_qual: out    vl_logic;
        lsc_prog_cipher_key1_qual: out    vl_logic;
        lsc_prog_pubkey0_qual: out    vl_logic;
        lsc_prog_pubkey1_qual: out    vl_logic;
        lsc_prog_pubkey2_qual: out    vl_logic;
        lsc_prog_pubkey3_qual: out    vl_logic;
        lsc_prog_feature_qual: out    vl_logic;
        lsc_prog_feabits_qual: out    vl_logic;
        lsc_prog_trim0_qual: out    vl_logic;
        lsc_prog_trim1_qual: out    vl_logic;
        lsc_prog_pes_qual: out    vl_logic;
        lsc_prog_mes_qual: out    vl_logic;
        lsc_prog_usec_qual: out    vl_logic;
        lsc_prog_csec_qual: out    vl_logic;
        lsc_prog_uds_qual: out    vl_logic;
        lsc_read_authmode_qual: out    vl_logic;
        lsc_read_aesfea_qual: out    vl_logic;
        lsc_read_password_qual: out    vl_logic;
        lsc_read_cipher_key0_qual: out    vl_logic;
        lsc_read_cipher_key1_qual: out    vl_logic;
        lsc_read_pubkey0_qual: out    vl_logic;
        lsc_read_pubkey1_qual: out    vl_logic;
        lsc_read_pubkey2_qual: out    vl_logic;
        lsc_read_pubkey3_qual: out    vl_logic;
        lsc_read_feature_qual: out    vl_logic;
        lsc_read_feabits_qual: out    vl_logic;
        lsc_read_trim0_qual: out    vl_logic;
        lsc_read_trim1_qual: out    vl_logic;
        lsc_read_pes_qual: out    vl_logic;
        lsc_read_mes_qual: out    vl_logic;
        lsc_read_usec_qual: out    vl_logic;
        lsc_read_csec_qual: out    vl_logic;
        mfg_mdata_qual  : out    vl_logic;
        mfg_mtrim_qual  : out    vl_logic;
        cmd_read_exec_buf: out    vl_logic;
        cmd_read_cfg_reg: out    vl_logic;
        cmd_prog_cfg_reg: out    vl_logic;
        bse_prog_incr_cqual: out    vl_logic;
        lsc_i2ci_crbr_wt_qual: out    vl_logic;
        lsc_i2ci_txdr_wt_qual: out    vl_logic;
        lsc_i2ci_rxdr_rd_qual: out    vl_logic;
        lsc_i2ci_sr_rd_qual: out    vl_logic;
        lsc_read_i2c_qual: out    vl_logic;
        lsc_auth_ctrl_cqual: out    vl_logic;
        fl_prog_pubkey0_qual: out    vl_logic;
        fl_prog_pubkey1_qual: out    vl_logic;
        fl_prog_pubkey2_qual: out    vl_logic;
        fl_prog_pubkey3_qual: out    vl_logic;
        cmd_altsec_sram : out    vl_logic;
        cmd_altsec_cfg0 : out    vl_logic;
        cmd_altsec_cfg1 : out    vl_logic;
        cmd_altsec_ufm0 : out    vl_logic;
        cmd_altsec_ufm1 : out    vl_logic;
        cmd_altsec_ufm2 : out    vl_logic;
        cmd_altsec_ufm3 : out    vl_logic;
        cmd_altsec_trim : out    vl_logic;
        cmd_altsec_fea  : out    vl_logic;
        cmd_altsec_pubkey: out    vl_logic;
        cmd_altsec_aeskey: out    vl_logic;
        cmd_altsec_usec : out    vl_logic;
        cmd_altsec_csec : out    vl_logic;
        cmd_altsec_jtag : out    vl_logic;
        cmd_altsec_sspi : out    vl_logic;
        cmd_altsec_si2c : out    vl_logic;
        cmd_altsec_bspi : out    vl_logic;
        cmd_altsec_bi2c : out    vl_logic;
        sector_erase_pre: out    vl_logic_vector(11 downto 0);
        stat_sec_code   : out    vl_logic_vector(3 downto 0);
        stat_sec_bits   : out    vl_logic_vector(3 downto 0);
        stat_read_en    : out    vl_logic;
        stat_write_en   : out    vl_logic;
        stat_erase_en   : out    vl_logic;
        qualFail        : out    vl_logic;
        scanen          : in     vl_logic;
        sram_sec_prog   : in     vl_logic;
        sram_sec_read   : in     vl_logic;
        sd_sec_read_sram: in     vl_logic;
        sd_sec_erase_sram: in     vl_logic;
        sd_sec_hlock_sram: in     vl_logic;
        sd_sec_read_cfg0: in     vl_logic;
        sd_sec_prog_cfg0: in     vl_logic;
        sd_sec_erase_cfg0: in     vl_logic;
        sd_sec_hlock_cfg0: in     vl_logic;
        sd_sec_read_cfg1: in     vl_logic;
        sd_sec_prog_cfg1: in     vl_logic;
        sd_sec_erase_cfg1: in     vl_logic;
        sd_sec_hlock_cfg1: in     vl_logic;
        sd_sec_read_ufm0: in     vl_logic;
        sd_sec_prog_ufm0: in     vl_logic;
        sd_sec_erase_ufm0: in     vl_logic;
        sd_sec_hlock_ufm0: in     vl_logic;
        sd_sec_read_ufm1: in     vl_logic;
        sd_sec_prog_ufm1: in     vl_logic;
        sd_sec_erase_ufm1: in     vl_logic;
        sd_sec_hlock_ufm1: in     vl_logic;
        sd_sec_read_ufm2: in     vl_logic;
        sd_sec_prog_ufm2: in     vl_logic;
        sd_sec_erase_ufm2: in     vl_logic;
        sd_sec_hlock_ufm2: in     vl_logic;
        sd_sec_read_ufm3: in     vl_logic;
        sd_sec_prog_ufm3: in     vl_logic;
        sd_sec_erase_ufm3: in     vl_logic;
        sd_sec_hlock_ufm3: in     vl_logic;
        sd_sec_read_trim: in     vl_logic;
        sd_sec_prog_trim: in     vl_logic;
        sd_sec_erase_trim: in     vl_logic;
        sd_sec_hlock_trim: in     vl_logic;
        sd_sec_read_fea : in     vl_logic;
        sd_sec_prog_fea : in     vl_logic;
        sd_sec_erase_fea: in     vl_logic;
        sd_sec_hlock_fea: in     vl_logic;
        sd_sec_read_pubkey: in     vl_logic;
        sd_sec_prog_pubkey: in     vl_logic;
        sd_sec_erase_pubkey: in     vl_logic;
        sd_sec_hlock_pubkey: in     vl_logic;
        sd_sec_read_aeskey: in     vl_logic;
        sd_sec_prog_aeskey: in     vl_logic;
        sd_sec_erase_aeskey: in     vl_logic;
        sd_sec_hlock_aeskey: in     vl_logic;
        sd_sec_read_usec: in     vl_logic;
        sd_sec_prog_usec: in     vl_logic;
        sd_sec_erase_usec: in     vl_logic;
        sd_sec_hlock_usec: in     vl_logic;
        sd_sec_read_csec: in     vl_logic;
        sd_sec_prog_csec: in     vl_logic;
        sd_sec_erase_csec: in     vl_logic;
        sd_sec_hlock_csec: in     vl_logic;
        sd_sec_hlock_jtag: in     vl_logic;
        sd_sec_hlock_sspi: in     vl_logic;
        sd_sec_hlock_si2c: in     vl_logic;
        sd_sec_hlock_bspi: in     vl_logic;
        sd_sec_hlock_bi2c: in     vl_logic;
        sd_pwd_mismatch : in     vl_logic;
        sd_pwd_all      : in     vl_logic;
        sd_pwd_ufm      : in     vl_logic;
        sd_secplus_cfg0 : in     vl_logic;
        sd_secplus_cfg1 : in     vl_logic;
        sd_dec_only     : in     vl_logic;
        sd_auth_en      : in     vl_logic_vector(1 downto 0);
        sd_authdone_cfg0: in     vl_logic;
        sd_authdone_cfg1: in     vl_logic;
        bse_active      : in     vl_logic;
        fl_busy_sdm     : in     vl_logic;
        mstr_busy_bse   : in     vl_logic;
        njbse_rxdec     : in     vl_logic;
        mfg_margin      : in     vl_logic;
        p_mspi_all      : in     vl_logic;
        isc_exec_d      : in     vl_logic;
        isc_exec_e      : in     vl_logic;
        isc_exec_c      : in     vl_logic;
        dryrun_inp      : in     vl_logic;
        spi_flash_check_inp: in     vl_logic;
        cfg_sed_en      : in     vl_logic;
        access_sram     : in     vl_logic;
        access_flash    : in     vl_logic;
        access_tag      : in     vl_logic;
        current_sector  : in     vl_logic_vector(11 downto 0);
        sector_dat      : in     vl_logic_vector(15 downto 0);
        isc_data_shift_iq: in     vl_logic;
        isc_addr_shift_iq: in     vl_logic;
        verify_id_iq    : in     vl_logic;
        read_temp_iq    : in     vl_logic;
        lsc_device_ctrl_iq: in     vl_logic;
        prog_dryrun_addr_iq: in     vl_logic;
        lsc_shift_password_iq: in     vl_logic;
        lsc_bitstream_burst_iq: in     vl_logic;
        lsc_i2ci_crbr_wt_iq: in     vl_logic;
        lsc_i2ci_txdr_wt_iq: in     vl_logic;
        lsc_i2ci_rxdr_rd_iq: in     vl_logic;
        lsc_i2ci_sr_rd_iq: in     vl_logic;
        lsc_read_pes_mq : in     vl_logic;
        lsc_prog_ctrl0_iq: in     vl_logic;
        lsc_read_ctrl0_iq: in     vl_logic;
        lsc_prog_ctrl1_iq: in     vl_logic;
        lsc_read_ctrl1_iq: in     vl_logic;
        lsc_reset_crc_iq: in     vl_logic;
        lsc_read_crc_iq : in     vl_logic;
        lsc_write_comp_dic_iq: in     vl_logic;
        lsc_read_comp_dic_mq: in     vl_logic;
        sf_prog_ucode_iq: in     vl_logic;
        sf_program_iq   : in     vl_logic;
        sf_read_iq      : in     vl_logic;
        sf_erase_iq     : in     vl_logic;
        sf_prog_done_iq : in     vl_logic;
        sf_erase_done_iq: in     vl_logic;
        sf_prog_sec_iq  : in     vl_logic;
        sf_init_addr_iq : in     vl_logic;
        sf_write_addr_iq: in     vl_logic;
        sf_prog_incr_rti_iq: in     vl_logic;
        sf_prog_incr_enc_iq: in     vl_logic;
        sf_prog_incr_cmp_iq: in     vl_logic;
        sf_prog_incr_cne_iq: in     vl_logic;
        sf_vfy_incr_rti_iq: in     vl_logic;
        sf_prog_sed_crc_iq: in     vl_logic;
        sf_read_sed_crc_iq: in     vl_logic;
        sf_write_bus_addr_iq: in     vl_logic;
        sf_pcs_write_iq : in     vl_logic;
        sf_pcs_read_iq  : in     vl_logic;
        sf_ebr_write_iq : in     vl_logic;
        sf_ebr_read_iq  : in     vl_logic;
        fl_erase_iq     : in     vl_logic;
        fl_prog_done_iq : in     vl_logic;
        fl_prog_sec_iq  : in     vl_logic;
        fl_prog_secplus_iq: in     vl_logic;
        fl_prog_ucode_iq: in     vl_logic;
        fl_init_addr_iq : in     vl_logic;
        fl_write_addr_iq: in     vl_logic;
        fl_prog_incr_nv_iq: in     vl_logic;
        fl_read_incr_nv_iq: in     vl_logic;
        fl_prog_password_iq: in     vl_logic;
        fl_read_password_iq: in     vl_logic;
        fl_prog_cipher_key0_iq: in     vl_logic;
        fl_read_cipher_key0_iq: in     vl_logic;
        fl_prog_cipher_key1_iq: in     vl_logic;
        fl_read_cipher_key1_iq: in     vl_logic;
        fl_prog_feature_iq: in     vl_logic;
        fl_read_feature_iq: in     vl_logic;
        fl_prog_feabits_iq: in     vl_logic;
        fl_read_feabits_iq: in     vl_logic;
        fl_init_addr_ufm_iq: in     vl_logic;
        fl_prog_tag_iq  : in     vl_logic;
        fl_erase_tag_iq : in     vl_logic;
        fl_read_tag_iq  : in     vl_logic;
        fl_prog_pes_mq  : in     vl_logic;
        fl_prog_trim0_mq: in     vl_logic;
        fl_prog_trim1_mq: in     vl_logic;
        fl_prog_mes_mq  : in     vl_logic;
        fl_prog_hes_mq  : in     vl_logic;
        fl_read_trim0_mq: in     vl_logic;
        fl_read_trim1_mq: in     vl_logic;
        fl_read_mes_mq  : in     vl_logic;
        fl_read_hes_mq  : in     vl_logic;
        fl_prog_csec_iq : in     vl_logic;
        fl_read_csec_iq : in     vl_logic;
        fl_prog_usec_iq : in     vl_logic;
        fl_read_usec_iq : in     vl_logic;
        fl_prog_authdone_iq: in     vl_logic;
        fl_prog_authmode_iq: in     vl_logic;
        fl_prog_aesfea_iq: in     vl_logic;
        fl_read_authmode_iq: in     vl_logic;
        fl_read_aesfea_iq: in     vl_logic;
        mfg_en          : in     vl_logic;
        mfg_mtest_mq    : in     vl_logic;
        mfg_mtrim_mq    : in     vl_logic;
        mfg_mdata_mq    : in     vl_logic;
        isc_data_shift_cq: in     vl_logic;
        isc_addr_shift_cq: in     vl_logic;
        verify_id_cq    : in     vl_logic;
        read_temp_cq    : in     vl_logic;
        lsc_device_ctrl_cq: in     vl_logic;
        prog_dryrun_addr_cq: in     vl_logic;
        lsc_shift_password_cq: in     vl_logic;
        lsc_bitstream_burst_cq: in     vl_logic;
        lsc_read_pes_cq : in     vl_logic;
        lsc_prog_ctrl0_cq: in     vl_logic;
        lsc_read_ctrl0_cq: in     vl_logic;
        lsc_prog_ctrl1_cq: in     vl_logic;
        lsc_read_ctrl1_cq: in     vl_logic;
        lsc_reset_crc_cq: in     vl_logic;
        lsc_read_crc_cq : in     vl_logic;
        lsc_write_comp_dic_cq: in     vl_logic;
        sf_prog_ucode_cq: in     vl_logic;
        sf_program_cq   : in     vl_logic;
        sf_read_cq      : in     vl_logic;
        sf_erase_cq     : in     vl_logic;
        sf_prog_done_cq : in     vl_logic;
        sf_erase_done_cq: in     vl_logic;
        sf_prog_sec_cq  : in     vl_logic;
        sf_init_addr_cq : in     vl_logic;
        sf_write_addr_cq: in     vl_logic;
        sf_prog_incr_rti_cq: in     vl_logic;
        sf_prog_incr_enc_cq: in     vl_logic;
        sf_prog_incr_cmp_cq: in     vl_logic;
        sf_prog_incr_cne_cq: in     vl_logic;
        sf_vfy_incr_rti_cq: in     vl_logic;
        sf_prog_sed_crc_cq: in     vl_logic;
        sf_read_sed_crc_cq: in     vl_logic;
        sf_write_bus_addr_cq: in     vl_logic;
        sf_pcs_write_cq : in     vl_logic;
        sf_pcs_read_cq  : in     vl_logic;
        sf_ebr_write_cq : in     vl_logic;
        sf_ebr_read_cq  : in     vl_logic;
        fl_erase_cq     : in     vl_logic;
        fl_prog_done_cq : in     vl_logic;
        fl_prog_sec_cq  : in     vl_logic;
        fl_prog_secplus_cq: in     vl_logic;
        fl_prog_ucode_cq: in     vl_logic;
        fl_init_addr_cq : in     vl_logic;
        fl_write_addr_cq: in     vl_logic;
        fl_prog_incr_nv_cq: in     vl_logic;
        fl_read_incr_nv_cq: in     vl_logic;
        fl_prog_password_cq: in     vl_logic;
        fl_read_password_cq: in     vl_logic;
        fl_prog_cipher_key0_cq: in     vl_logic;
        fl_read_cipher_key0_cq: in     vl_logic;
        fl_prog_cipher_key1_cq: in     vl_logic;
        fl_read_cipher_key1_cq: in     vl_logic;
        fl_prog_feature_cq: in     vl_logic;
        fl_read_feature_cq: in     vl_logic;
        fl_prog_feabits_cq: in     vl_logic;
        fl_read_feabits_cq: in     vl_logic;
        fl_init_addr_ufm_cq: in     vl_logic;
        fl_prog_tag_cq  : in     vl_logic;
        fl_erase_tag_cq : in     vl_logic;
        fl_read_tag_cq  : in     vl_logic;
        fl_prog_csec_cq : in     vl_logic;
        fl_read_csec_cq : in     vl_logic;
        fl_prog_usec_cq : in     vl_logic;
        fl_read_usec_cq : in     vl_logic;
        fl_prog_authdone_cq: in     vl_logic;
        fl_prog_authmode_cq: in     vl_logic;
        fl_prog_aesfea_cq: in     vl_logic;
        fl_read_authmode_cq: in     vl_logic;
        fl_read_aesfea_cq: in     vl_logic;
        lsc_jump_cq     : in     vl_logic;
        lsc_chip_select_cq: in     vl_logic;
        lsc_flow_through_cq: in     vl_logic;
        bypass_cq       : in     vl_logic;
        sed_init_addr_cq: in     vl_logic;
        sed_write_addr_cq: in     vl_logic;
        sed_prog_incr_rti_cq: in     vl_logic;
        sed_prog_incr_cmp_cq: in     vl_logic;
        sed_prog_sed_crc_cq: in     vl_logic;
        sed_prog_ctrl0_cq: in     vl_logic;
        sed_prog_ctrl1_cq: in     vl_logic;
        sed_write_comp_dic_cq: in     vl_logic;
        lsc_i2ci_crbr_wt_cq: in     vl_logic;
        lsc_i2ci_txdr_wt_cq: in     vl_logic;
        lsc_i2ci_rxdr_rd_cq: in     vl_logic;
        lsc_i2ci_sr_rd_cq: in     vl_logic;
        lsc_alter_sec_cq: in     vl_logic;
        lsc_alter_sram_sec_cq: in     vl_logic;
        lsc_alter_port_sec_cq: in     vl_logic;
        lsc_prog_uds_cq : in     vl_logic;
        uds_trn_blank   : in     vl_logic;
        hse_trn_valid   : in     vl_logic;
        lsc_auth_ctrl_cq: in     vl_logic;
        fl_prog_pubkey0_cq: in     vl_logic;
        fl_read_pubkey0_cq: in     vl_logic;
        fl_prog_pubkey1_cq: in     vl_logic;
        fl_read_pubkey1_cq: in     vl_logic;
        fl_prog_pubkey2_cq: in     vl_logic;
        fl_read_pubkey2_cq: in     vl_logic;
        fl_prog_pubkey3_cq: in     vl_logic;
        fl_read_pubkey3_cq: in     vl_logic;
        fl_prog_pubkey0_iq: in     vl_logic;
        fl_read_pubkey0_iq: in     vl_logic;
        fl_prog_pubkey1_iq: in     vl_logic;
        fl_read_pubkey1_iq: in     vl_logic;
        fl_prog_pubkey2_iq: in     vl_logic;
        fl_read_pubkey2_iq: in     vl_logic;
        fl_prog_pubkey3_iq: in     vl_logic;
        fl_read_pubkey3_iq: in     vl_logic;
        wbc_active      : in     vl_logic
    );
end cfg_qual;
