library verilog;
use verilog.vl_types.all;
entity SYSBUSA_sim is
    generic(
        SYSBUS_CONFIG_FILE: string  := "sysbuscfgfile.txt";
        BASE_ADDRESS    : string  := "0x3EF00";
        MPI_PARITY      : string  := "DISABLED";
        MPI_BUS_WIDTH   : integer := 8;
        SYS_CLK_SEL     : string  := "MPI";
        MPI_PRIORITY    : string  := "LOW";
        FPGA_PRIORITY   : string  := "LOW";
        MPI_RST         : string  := "DISABLED";
        MASTER_RST      : string  := "DISABLED";
        PARITY          : string  := "EVEN";
        MPI_SYNCMODE    : string  := "SYNC";
        MASTER_SYNCMODE : string  := "ASYNC";
        MASTER_AUTORETRY: string  := "ENABLED";
        SLAVE_SYNCMODE  : string  := "ASYNC";
        INTERRUPT_VECTOR1: integer := 0;
        INTERRUPT_VECTOR2: integer := 0;
        INTERRUPT_VECTOR3: integer := 0;
        INTERRUPT_VECTOR4: integer := 0;
        INTERRUPT_VECTOR5: integer := 0;
        INTERRUPT_VECTOR6: integer := 0;
        WS_TIME_INDEX   : integer := 4;
        GRANT_TIME_INDEX: integer := 0
    );
    port(
        CS0_N           : in     vl_logic;
        CS1             : in     vl_logic;
        MPI_CLK         : in     vl_logic;
        MPI_WR_N        : in     vl_logic;
        MPI_STRB_N      : in     vl_logic;
        MPI_TSIZ_1      : in     vl_logic;
        MPI_TSIZ_0      : in     vl_logic;
        MPI_BURST       : in     vl_logic;
        MPI_BDIP        : in     vl_logic;
        MPI_ADDR_14     : in     vl_logic;
        MPI_ADDR_15     : in     vl_logic;
        MPI_ADDR_16     : in     vl_logic;
        MPI_ADDR_17     : in     vl_logic;
        MPI_ADDR_18     : in     vl_logic;
        MPI_ADDR_19     : in     vl_logic;
        MPI_ADDR_20     : in     vl_logic;
        MPI_ADDR_21     : in     vl_logic;
        MPI_ADDR_22     : in     vl_logic;
        MPI_ADDR_23     : in     vl_logic;
        MPI_ADDR_24     : in     vl_logic;
        MPI_ADDR_25     : in     vl_logic;
        MPI_ADDR_26     : in     vl_logic;
        MPI_ADDR_27     : in     vl_logic;
        MPI_ADDR_28     : in     vl_logic;
        MPI_ADDR_29     : in     vl_logic;
        MPI_ADDR_30     : in     vl_logic;
        MPI_ADDR_31     : in     vl_logic;
        MPI_WR_DATA_31  : in     vl_logic;
        MPI_WR_DATA_30  : in     vl_logic;
        MPI_WR_DATA_29  : in     vl_logic;
        MPI_WR_DATA_28  : in     vl_logic;
        MPI_WR_DATA_27  : in     vl_logic;
        MPI_WR_DATA_26  : in     vl_logic;
        MPI_WR_DATA_25  : in     vl_logic;
        MPI_WR_DATA_24  : in     vl_logic;
        MPI_WR_DATA_23  : in     vl_logic;
        MPI_WR_DATA_22  : in     vl_logic;
        MPI_WR_DATA_21  : in     vl_logic;
        MPI_WR_DATA_20  : in     vl_logic;
        MPI_WR_DATA_19  : in     vl_logic;
        MPI_WR_DATA_18  : in     vl_logic;
        MPI_WR_DATA_17  : in     vl_logic;
        MPI_WR_DATA_16  : in     vl_logic;
        MPI_WR_DATA_15  : in     vl_logic;
        MPI_WR_DATA_14  : in     vl_logic;
        MPI_WR_DATA_13  : in     vl_logic;
        MPI_WR_DATA_12  : in     vl_logic;
        MPI_WR_DATA_11  : in     vl_logic;
        MPI_WR_DATA_10  : in     vl_logic;
        MPI_WR_DATA_9   : in     vl_logic;
        MPI_WR_DATA_8   : in     vl_logic;
        MPI_WR_DATA_7   : in     vl_logic;
        MPI_WR_DATA_6   : in     vl_logic;
        MPI_WR_DATA_5   : in     vl_logic;
        MPI_WR_DATA_4   : in     vl_logic;
        MPI_WR_DATA_3   : in     vl_logic;
        MPI_WR_DATA_2   : in     vl_logic;
        MPI_WR_DATA_1   : in     vl_logic;
        MPI_WR_DATA_0   : in     vl_logic;
        MPI_WR_PARITY_3 : in     vl_logic;
        MPI_WR_PARITY_2 : in     vl_logic;
        MPI_WR_PARITY_1 : in     vl_logic;
        MPI_WR_PARITY_0 : in     vl_logic;
        MPI_RST_N       : in     vl_logic;
        SYS_RST_N       : in     vl_logic;
        USR_CLK         : in     vl_logic;
        USER_IRQ_IN     : in     vl_logic;
        MPI_TA          : out    vl_logic;
        MPI_RETRY       : out    vl_logic;
        MPI_TEA         : out    vl_logic;
        MPI_RD_DATA_31  : out    vl_logic;
        MPI_RD_DATA_30  : out    vl_logic;
        MPI_RD_DATA_29  : out    vl_logic;
        MPI_RD_DATA_28  : out    vl_logic;
        MPI_RD_DATA_27  : out    vl_logic;
        MPI_RD_DATA_26  : out    vl_logic;
        MPI_RD_DATA_25  : out    vl_logic;
        MPI_RD_DATA_24  : out    vl_logic;
        MPI_RD_DATA_23  : out    vl_logic;
        MPI_RD_DATA_22  : out    vl_logic;
        MPI_RD_DATA_21  : out    vl_logic;
        MPI_RD_DATA_20  : out    vl_logic;
        MPI_RD_DATA_19  : out    vl_logic;
        MPI_RD_DATA_18  : out    vl_logic;
        MPI_RD_DATA_17  : out    vl_logic;
        MPI_RD_DATA_16  : out    vl_logic;
        MPI_RD_DATA_15  : out    vl_logic;
        MPI_RD_DATA_14  : out    vl_logic;
        MPI_RD_DATA_13  : out    vl_logic;
        MPI_RD_DATA_12  : out    vl_logic;
        MPI_RD_DATA_11  : out    vl_logic;
        MPI_RD_DATA_10  : out    vl_logic;
        MPI_RD_DATA_9   : out    vl_logic;
        MPI_RD_DATA_8   : out    vl_logic;
        MPI_RD_DATA_7   : out    vl_logic;
        MPI_RD_DATA_6   : out    vl_logic;
        MPI_RD_DATA_5   : out    vl_logic;
        MPI_RD_DATA_4   : out    vl_logic;
        MPI_RD_DATA_3   : out    vl_logic;
        MPI_RD_DATA_2   : out    vl_logic;
        MPI_RD_DATA_1   : out    vl_logic;
        MPI_RD_DATA_0   : out    vl_logic;
        PD2_0_TS        : out    vl_logic;
        PD7_3_TS        : out    vl_logic;
        PD15_8_TS       : out    vl_logic;
        PD31_16_TS      : out    vl_logic;
        MPI_RD_PARITY_3 : out    vl_logic;
        MPI_RD_PARITY_2 : out    vl_logic;
        MPI_RD_PARITY_1 : out    vl_logic;
        MPI_RD_PARITY_0 : out    vl_logic;
        MPI_DP_TS_0     : out    vl_logic;
        MPI_DP_TS_1     : out    vl_logic;
        MPI_DP_TS_2     : out    vl_logic;
        MPI_IRQ_N       : out    vl_logic;
        MPI_CNTL_TS     : out    vl_logic;
        USER_IRQ_OUT    : out    vl_logic;
        HCLK_CIB        : out    vl_logic;
        SMI_RDATA_63    : in     vl_logic;
        SMI_RDATA_62    : in     vl_logic;
        SMI_RDATA_61    : in     vl_logic;
        SMI_RDATA_60    : in     vl_logic;
        SMI_RDATA_59    : in     vl_logic;
        SMI_RDATA_58    : in     vl_logic;
        SMI_RDATA_57    : in     vl_logic;
        SMI_RDATA_56    : in     vl_logic;
        SMI_RDATA_55    : in     vl_logic;
        SMI_RDATA_54    : in     vl_logic;
        SMI_RDATA_53    : in     vl_logic;
        SMI_RDATA_52    : in     vl_logic;
        SMI_RDATA_51    : in     vl_logic;
        SMI_RDATA_50    : in     vl_logic;
        SMI_RDATA_49    : in     vl_logic;
        SMI_RDATA_48    : in     vl_logic;
        SMI_RDATA_47    : in     vl_logic;
        SMI_RDATA_46    : in     vl_logic;
        SMI_RDATA_45    : in     vl_logic;
        SMI_RDATA_44    : in     vl_logic;
        SMI_RDATA_43    : in     vl_logic;
        SMI_RDATA_42    : in     vl_logic;
        SMI_RDATA_41    : in     vl_logic;
        SMI_RDATA_40    : in     vl_logic;
        SMI_RDATA_39    : in     vl_logic;
        SMI_RDATA_38    : in     vl_logic;
        SMI_RDATA_37    : in     vl_logic;
        SMI_RDATA_36    : in     vl_logic;
        SMI_RDATA_35    : in     vl_logic;
        SMI_RDATA_34    : in     vl_logic;
        SMI_RDATA_33    : in     vl_logic;
        SMI_RDATA_32    : in     vl_logic;
        SMI_RDATA_31    : in     vl_logic;
        SMI_RDATA_30    : in     vl_logic;
        SMI_RDATA_29    : in     vl_logic;
        SMI_RDATA_28    : in     vl_logic;
        SMI_RDATA_27    : in     vl_logic;
        SMI_RDATA_26    : in     vl_logic;
        SMI_RDATA_25    : in     vl_logic;
        SMI_RDATA_24    : in     vl_logic;
        SMI_RDATA_23    : in     vl_logic;
        SMI_RDATA_22    : in     vl_logic;
        SMI_RDATA_21    : in     vl_logic;
        SMI_RDATA_20    : in     vl_logic;
        SMI_RDATA_19    : in     vl_logic;
        SMI_RDATA_18    : in     vl_logic;
        SMI_RDATA_17    : in     vl_logic;
        SMI_RDATA_16    : in     vl_logic;
        SMI_RDATA_15    : in     vl_logic;
        SMI_RDATA_14    : in     vl_logic;
        SMI_RDATA_13    : in     vl_logic;
        SMI_RDATA_12    : in     vl_logic;
        SMI_RDATA_11    : in     vl_logic;
        SMI_RDATA_10    : in     vl_logic;
        SMI_RDATA_9     : in     vl_logic;
        SMI_RDATA_8     : in     vl_logic;
        SMI_RDATA_7     : in     vl_logic;
        SMI_RDATA_6     : in     vl_logic;
        SMI_RDATA_5     : in     vl_logic;
        SMI_RDATA_4     : in     vl_logic;
        SMI_RDATA_3     : in     vl_logic;
        SMI_RDATA_2     : in     vl_logic;
        SMI_RDATA_1     : in     vl_logic;
        SMI_RDATA_0     : in     vl_logic;
        SMI_ADDR_9      : out    vl_logic;
        SMI_ADDR_8      : out    vl_logic;
        SMI_ADDR_7      : out    vl_logic;
        SMI_ADDR_6      : out    vl_logic;
        SMI_ADDR_5      : out    vl_logic;
        SMI_ADDR_4      : out    vl_logic;
        SMI_ADDR_3      : out    vl_logic;
        SMI_ADDR_2      : out    vl_logic;
        SMI_ADDR_1      : out    vl_logic;
        SMI_ADDR_0      : out    vl_logic;
        SMI_CLK         : out    vl_logic;
        SMI_RD          : out    vl_logic;
        SMI_RST_N       : out    vl_logic;
        SMI_WDATA       : out    vl_logic;
        SMI_WR          : out    vl_logic;
        FMADDR_0        : in     vl_logic;
        FMADDR_1        : in     vl_logic;
        FMADDR_2        : in     vl_logic;
        FMADDR_3        : in     vl_logic;
        FMADDR_4        : in     vl_logic;
        FMADDR_5        : in     vl_logic;
        FMADDR_6        : in     vl_logic;
        FMADDR_7        : in     vl_logic;
        FMADDR_8        : in     vl_logic;
        FMADDR_9        : in     vl_logic;
        FMADDR_10       : in     vl_logic;
        FMADDR_11       : in     vl_logic;
        FMADDR_12       : in     vl_logic;
        FMADDR_13       : in     vl_logic;
        FMADDR_14       : in     vl_logic;
        FMADDR_15       : in     vl_logic;
        FMADDR_16       : in     vl_logic;
        FMADDR_17       : in     vl_logic;
        FMWDATA_0       : in     vl_logic;
        FMWDATA_1       : in     vl_logic;
        FMWDATA_2       : in     vl_logic;
        FMWDATA_3       : in     vl_logic;
        FMWDATA_4       : in     vl_logic;
        FMWDATA_5       : in     vl_logic;
        FMWDATA_6       : in     vl_logic;
        FMWDATA_7       : in     vl_logic;
        FMWDATA_8       : in     vl_logic;
        FMWDATA_9       : in     vl_logic;
        FMWDATA_10      : in     vl_logic;
        FMWDATA_11      : in     vl_logic;
        FMWDATA_12      : in     vl_logic;
        FMWDATA_13      : in     vl_logic;
        FMWDATA_14      : in     vl_logic;
        FMWDATA_15      : in     vl_logic;
        FMWDATA_16      : in     vl_logic;
        FMWDATA_17      : in     vl_logic;
        FMWDATA_18      : in     vl_logic;
        FMWDATA_19      : in     vl_logic;
        FMWDATA_20      : in     vl_logic;
        FMWDATA_21      : in     vl_logic;
        FMWDATA_22      : in     vl_logic;
        FMWDATA_23      : in     vl_logic;
        FMWDATA_24      : in     vl_logic;
        FMWDATA_25      : in     vl_logic;
        FMWDATA_26      : in     vl_logic;
        FMWDATA_27      : in     vl_logic;
        FMWDATA_28      : in     vl_logic;
        FMWDATA_29      : in     vl_logic;
        FMWDATA_30      : in     vl_logic;
        FMWDATA_31      : in     vl_logic;
        FMWDATA_32      : in     vl_logic;
        FMWDATA_33      : in     vl_logic;
        FMWDATA_34      : in     vl_logic;
        FMWDATA_35      : in     vl_logic;
        FMCLK           : in     vl_logic;
        FMRESET_N       : in     vl_logic;
        FMWRN           : in     vl_logic;
        FMBURST         : in     vl_logic;
        FMRDY           : in     vl_logic;
        FMSIZE_0        : in     vl_logic;
        FMSIZE_1        : in     vl_logic;
        FMLOCK          : in     vl_logic;
        FMIRQ           : in     vl_logic;
        FMRDATA_0       : out    vl_logic;
        FMRDATA_1       : out    vl_logic;
        FMRDATA_2       : out    vl_logic;
        FMRDATA_3       : out    vl_logic;
        FMRDATA_4       : out    vl_logic;
        FMRDATA_5       : out    vl_logic;
        FMRDATA_6       : out    vl_logic;
        FMRDATA_7       : out    vl_logic;
        FMRDATA_8       : out    vl_logic;
        FMRDATA_9       : out    vl_logic;
        FMRDATA_10      : out    vl_logic;
        FMRDATA_11      : out    vl_logic;
        FMRDATA_12      : out    vl_logic;
        FMRDATA_13      : out    vl_logic;
        FMRDATA_14      : out    vl_logic;
        FMRDATA_15      : out    vl_logic;
        FMRDATA_16      : out    vl_logic;
        FMRDATA_17      : out    vl_logic;
        FMRDATA_18      : out    vl_logic;
        FMRDATA_19      : out    vl_logic;
        FMRDATA_20      : out    vl_logic;
        FMRDATA_21      : out    vl_logic;
        FMRDATA_22      : out    vl_logic;
        FMRDATA_23      : out    vl_logic;
        FMRDATA_24      : out    vl_logic;
        FMRDATA_25      : out    vl_logic;
        FMRDATA_26      : out    vl_logic;
        FMRDATA_27      : out    vl_logic;
        FMRDATA_28      : out    vl_logic;
        FMRDATA_29      : out    vl_logic;
        FMRDATA_30      : out    vl_logic;
        FMRDATA_31      : out    vl_logic;
        FMRDATA_32      : out    vl_logic;
        FMRDATA_33      : out    vl_logic;
        FMRDATA_34      : out    vl_logic;
        FMRDATA_35      : out    vl_logic;
        FMACK           : out    vl_logic;
        FMRETRY         : out    vl_logic;
        FMERR           : out    vl_logic;
        FSRDATA_0       : in     vl_logic;
        FSRDATA_1       : in     vl_logic;
        FSRDATA_2       : in     vl_logic;
        FSRDATA_3       : in     vl_logic;
        FSRDATA_4       : in     vl_logic;
        FSRDATA_5       : in     vl_logic;
        FSRDATA_6       : in     vl_logic;
        FSRDATA_7       : in     vl_logic;
        FSRDATA_8       : in     vl_logic;
        FSRDATA_9       : in     vl_logic;
        FSRDATA_10      : in     vl_logic;
        FSRDATA_11      : in     vl_logic;
        FSRDATA_12      : in     vl_logic;
        FSRDATA_13      : in     vl_logic;
        FSRDATA_14      : in     vl_logic;
        FSRDATA_15      : in     vl_logic;
        FSRDATA_16      : in     vl_logic;
        FSRDATA_17      : in     vl_logic;
        FSRDATA_18      : in     vl_logic;
        FSRDATA_19      : in     vl_logic;
        FSRDATA_20      : in     vl_logic;
        FSRDATA_21      : in     vl_logic;
        FSRDATA_22      : in     vl_logic;
        FSRDATA_23      : in     vl_logic;
        FSRDATA_24      : in     vl_logic;
        FSRDATA_25      : in     vl_logic;
        FSRDATA_26      : in     vl_logic;
        FSRDATA_27      : in     vl_logic;
        FSRDATA_28      : in     vl_logic;
        FSRDATA_29      : in     vl_logic;
        FSRDATA_30      : in     vl_logic;
        FSRDATA_31      : in     vl_logic;
        FSRDATA_32      : in     vl_logic;
        FSRDATA_33      : in     vl_logic;
        FSRDATA_34      : in     vl_logic;
        FSRDATA_35      : in     vl_logic;
        FSCLK           : in     vl_logic;
        FSRESET_N       : in     vl_logic;
        FSACK           : in     vl_logic;
        FSRETRY         : in     vl_logic;
        FSERR           : in     vl_logic;
        FSIRQ           : in     vl_logic;
        FSWDATA_0       : out    vl_logic;
        FSWDATA_1       : out    vl_logic;
        FSWDATA_2       : out    vl_logic;
        FSWDATA_3       : out    vl_logic;
        FSWDATA_4       : out    vl_logic;
        FSWDATA_5       : out    vl_logic;
        FSWDATA_6       : out    vl_logic;
        FSWDATA_7       : out    vl_logic;
        FSWDATA_8       : out    vl_logic;
        FSWDATA_9       : out    vl_logic;
        FSWDATA_10      : out    vl_logic;
        FSWDATA_11      : out    vl_logic;
        FSWDATA_12      : out    vl_logic;
        FSWDATA_13      : out    vl_logic;
        FSWDATA_14      : out    vl_logic;
        FSWDATA_15      : out    vl_logic;
        FSWDATA_16      : out    vl_logic;
        FSWDATA_17      : out    vl_logic;
        FSWDATA_18      : out    vl_logic;
        FSWDATA_19      : out    vl_logic;
        FSWDATA_20      : out    vl_logic;
        FSWDATA_21      : out    vl_logic;
        FSWDATA_22      : out    vl_logic;
        FSWDATA_23      : out    vl_logic;
        FSWDATA_24      : out    vl_logic;
        FSWDATA_25      : out    vl_logic;
        FSWDATA_26      : out    vl_logic;
        FSWDATA_27      : out    vl_logic;
        FSWDATA_28      : out    vl_logic;
        FSWDATA_29      : out    vl_logic;
        FSWDATA_30      : out    vl_logic;
        FSWDATA_31      : out    vl_logic;
        FSWDATA_32      : out    vl_logic;
        FSWDATA_33      : out    vl_logic;
        FSWDATA_34      : out    vl_logic;
        FSWDATA_35      : out    vl_logic;
        FSADDR_0        : out    vl_logic;
        FSADDR_1        : out    vl_logic;
        FSADDR_2        : out    vl_logic;
        FSADDR_3        : out    vl_logic;
        FSADDR_4        : out    vl_logic;
        FSADDR_5        : out    vl_logic;
        FSADDR_6        : out    vl_logic;
        FSADDR_7        : out    vl_logic;
        FSADDR_8        : out    vl_logic;
        FSADDR_9        : out    vl_logic;
        FSADDR_10       : out    vl_logic;
        FSADDR_11       : out    vl_logic;
        FSADDR_12       : out    vl_logic;
        FSADDR_13       : out    vl_logic;
        FSADDR_14       : out    vl_logic;
        FSADDR_15       : out    vl_logic;
        FSADDR_16       : out    vl_logic;
        FSADDR_17       : out    vl_logic;
        FSRDY           : out    vl_logic;
        FSWRN           : out    vl_logic;
        FSSIZE_0        : out    vl_logic;
        FSSIZE_1        : out    vl_logic;
        HADDR_LASBM_17  : in     vl_logic;
        HADDR_LASBM_16  : in     vl_logic;
        HADDR_LASBM_15  : in     vl_logic;
        HADDR_LASBM_14  : in     vl_logic;
        HADDR_LASBM_13  : in     vl_logic;
        HADDR_LASBM_12  : in     vl_logic;
        HADDR_LASBM_11  : in     vl_logic;
        HADDR_LASBM_10  : in     vl_logic;
        HADDR_LASBM_9   : in     vl_logic;
        HADDR_LASBM_8   : in     vl_logic;
        HADDR_LASBM_7   : in     vl_logic;
        HADDR_LASBM_6   : in     vl_logic;
        HADDR_LASBM_5   : in     vl_logic;
        HADDR_LASBM_4   : in     vl_logic;
        HADDR_LASBM_3   : in     vl_logic;
        HADDR_LASBM_2   : in     vl_logic;
        HADDR_LASBM_1   : in     vl_logic;
        HADDR_LASBM_0   : in     vl_logic;
        HSIZE_LASBM_1   : in     vl_logic;
        HSIZE_LASBM_0   : in     vl_logic;
        HTRANS_LASBM_1  : in     vl_logic;
        HTRANS_LASBM_0  : in     vl_logic;
        HWDATA_LASBM_35 : in     vl_logic;
        HWDATA_LASBM_34 : in     vl_logic;
        HWDATA_LASBM_33 : in     vl_logic;
        HWDATA_LASBM_32 : in     vl_logic;
        HWDATA_LASBM_31 : in     vl_logic;
        HWDATA_LASBM_30 : in     vl_logic;
        HWDATA_LASBM_29 : in     vl_logic;
        HWDATA_LASBM_28 : in     vl_logic;
        HWDATA_LASBM_27 : in     vl_logic;
        HWDATA_LASBM_26 : in     vl_logic;
        HWDATA_LASBM_25 : in     vl_logic;
        HWDATA_LASBM_24 : in     vl_logic;
        HWDATA_LASBM_23 : in     vl_logic;
        HWDATA_LASBM_22 : in     vl_logic;
        HWDATA_LASBM_21 : in     vl_logic;
        HWDATA_LASBM_20 : in     vl_logic;
        HWDATA_LASBM_19 : in     vl_logic;
        HWDATA_LASBM_18 : in     vl_logic;
        HWDATA_LASBM_17 : in     vl_logic;
        HWDATA_LASBM_16 : in     vl_logic;
        HWDATA_LASBM_15 : in     vl_logic;
        HWDATA_LASBM_14 : in     vl_logic;
        HWDATA_LASBM_13 : in     vl_logic;
        HWDATA_LASBM_12 : in     vl_logic;
        HWDATA_LASBM_11 : in     vl_logic;
        HWDATA_LASBM_10 : in     vl_logic;
        HWDATA_LASBM_9  : in     vl_logic;
        HWDATA_LASBM_8  : in     vl_logic;
        HWDATA_LASBM_7  : in     vl_logic;
        HWDATA_LASBM_6  : in     vl_logic;
        HWDATA_LASBM_5  : in     vl_logic;
        HWDATA_LASBM_4  : in     vl_logic;
        HWDATA_LASBM_3  : in     vl_logic;
        HWDATA_LASBM_2  : in     vl_logic;
        HWDATA_LASBM_1  : in     vl_logic;
        HWDATA_LASBM_0  : in     vl_logic;
        HBURST_LASBM    : in     vl_logic;
        HWRITE_LASBM    : in     vl_logic;
        LASB_CLK        : in     vl_logic;
        LASB_GSR        : in     vl_logic;
        LASB_IRQ_MASTER : in     vl_logic;
        HRDATA_LASBM_35 : out    vl_logic;
        HRDATA_LASBM_34 : out    vl_logic;
        HRDATA_LASBM_33 : out    vl_logic;
        HRDATA_LASBM_32 : out    vl_logic;
        HRDATA_LASBM_31 : out    vl_logic;
        HRDATA_LASBM_30 : out    vl_logic;
        HRDATA_LASBM_29 : out    vl_logic;
        HRDATA_LASBM_28 : out    vl_logic;
        HRDATA_LASBM_27 : out    vl_logic;
        HRDATA_LASBM_26 : out    vl_logic;
        HRDATA_LASBM_25 : out    vl_logic;
        HRDATA_LASBM_24 : out    vl_logic;
        HRDATA_LASBM_23 : out    vl_logic;
        HRDATA_LASBM_22 : out    vl_logic;
        HRDATA_LASBM_21 : out    vl_logic;
        HRDATA_LASBM_20 : out    vl_logic;
        HRDATA_LASBM_19 : out    vl_logic;
        HRDATA_LASBM_18 : out    vl_logic;
        HRDATA_LASBM_17 : out    vl_logic;
        HRDATA_LASBM_16 : out    vl_logic;
        HRDATA_LASBM_15 : out    vl_logic;
        HRDATA_LASBM_14 : out    vl_logic;
        HRDATA_LASBM_13 : out    vl_logic;
        HRDATA_LASBM_12 : out    vl_logic;
        HRDATA_LASBM_11 : out    vl_logic;
        HRDATA_LASBM_10 : out    vl_logic;
        HRDATA_LASBM_9  : out    vl_logic;
        HRDATA_LASBM_8  : out    vl_logic;
        HRDATA_LASBM_7  : out    vl_logic;
        HRDATA_LASBM_6  : out    vl_logic;
        HRDATA_LASBM_5  : out    vl_logic;
        HRDATA_LASBM_4  : out    vl_logic;
        HRDATA_LASBM_3  : out    vl_logic;
        HRDATA_LASBM_2  : out    vl_logic;
        HRDATA_LASBM_1  : out    vl_logic;
        HRDATA_LASBM_0  : out    vl_logic;
        HRESP_LASBM_1   : out    vl_logic;
        HRESP_LASBM_0   : out    vl_logic;
        HCLK_LASB       : out    vl_logic;
        HREADY_LASB     : out    vl_logic;
        HRESET_N_LASB   : out    vl_logic;
        LASB_DONE       : out    vl_logic;
        LASB_GSR_N      : out    vl_logic;
        LASB_IRQ_OUT    : out    vl_logic;
        HADDR_RASBM_17  : in     vl_logic;
        HADDR_RASBM_16  : in     vl_logic;
        HADDR_RASBM_15  : in     vl_logic;
        HADDR_RASBM_14  : in     vl_logic;
        HADDR_RASBM_13  : in     vl_logic;
        HADDR_RASBM_12  : in     vl_logic;
        HADDR_RASBM_11  : in     vl_logic;
        HADDR_RASBM_10  : in     vl_logic;
        HADDR_RASBM_9   : in     vl_logic;
        HADDR_RASBM_8   : in     vl_logic;
        HADDR_RASBM_7   : in     vl_logic;
        HADDR_RASBM_6   : in     vl_logic;
        HADDR_RASBM_5   : in     vl_logic;
        HADDR_RASBM_4   : in     vl_logic;
        HADDR_RASBM_3   : in     vl_logic;
        HADDR_RASBM_2   : in     vl_logic;
        HADDR_RASBM_1   : in     vl_logic;
        HADDR_RASBM_0   : in     vl_logic;
        HSIZE_RASBM_1   : in     vl_logic;
        HSIZE_RASBM_0   : in     vl_logic;
        HTRANS_RASBM_1  : in     vl_logic;
        HTRANS_RASBM_0  : in     vl_logic;
        HWDATA_RASBM_35 : in     vl_logic;
        HWDATA_RASBM_34 : in     vl_logic;
        HWDATA_RASBM_33 : in     vl_logic;
        HWDATA_RASBM_32 : in     vl_logic;
        HWDATA_RASBM_31 : in     vl_logic;
        HWDATA_RASBM_30 : in     vl_logic;
        HWDATA_RASBM_29 : in     vl_logic;
        HWDATA_RASBM_28 : in     vl_logic;
        HWDATA_RASBM_27 : in     vl_logic;
        HWDATA_RASBM_26 : in     vl_logic;
        HWDATA_RASBM_25 : in     vl_logic;
        HWDATA_RASBM_24 : in     vl_logic;
        HWDATA_RASBM_23 : in     vl_logic;
        HWDATA_RASBM_22 : in     vl_logic;
        HWDATA_RASBM_21 : in     vl_logic;
        HWDATA_RASBM_20 : in     vl_logic;
        HWDATA_RASBM_19 : in     vl_logic;
        HWDATA_RASBM_18 : in     vl_logic;
        HWDATA_RASBM_17 : in     vl_logic;
        HWDATA_RASBM_16 : in     vl_logic;
        HWDATA_RASBM_15 : in     vl_logic;
        HWDATA_RASBM_14 : in     vl_logic;
        HWDATA_RASBM_13 : in     vl_logic;
        HWDATA_RASBM_12 : in     vl_logic;
        HWDATA_RASBM_11 : in     vl_logic;
        HWDATA_RASBM_10 : in     vl_logic;
        HWDATA_RASBM_9  : in     vl_logic;
        HWDATA_RASBM_8  : in     vl_logic;
        HWDATA_RASBM_7  : in     vl_logic;
        HWDATA_RASBM_6  : in     vl_logic;
        HWDATA_RASBM_5  : in     vl_logic;
        HWDATA_RASBM_4  : in     vl_logic;
        HWDATA_RASBM_3  : in     vl_logic;
        HWDATA_RASBM_2  : in     vl_logic;
        HWDATA_RASBM_1  : in     vl_logic;
        HWDATA_RASBM_0  : in     vl_logic;
        HBURST_RASBM    : in     vl_logic;
        HWRITE_RASBM    : in     vl_logic;
        RASB_CLK        : in     vl_logic;
        RASB_GSR        : in     vl_logic;
        RASB_IRQ_MASTER : in     vl_logic;
        HRDATA_RASBM_35 : out    vl_logic;
        HRDATA_RASBM_34 : out    vl_logic;
        HRDATA_RASBM_33 : out    vl_logic;
        HRDATA_RASBM_32 : out    vl_logic;
        HRDATA_RASBM_31 : out    vl_logic;
        HRDATA_RASBM_30 : out    vl_logic;
        HRDATA_RASBM_29 : out    vl_logic;
        HRDATA_RASBM_28 : out    vl_logic;
        HRDATA_RASBM_27 : out    vl_logic;
        HRDATA_RASBM_26 : out    vl_logic;
        HRDATA_RASBM_25 : out    vl_logic;
        HRDATA_RASBM_24 : out    vl_logic;
        HRDATA_RASBM_23 : out    vl_logic;
        HRDATA_RASBM_22 : out    vl_logic;
        HRDATA_RASBM_21 : out    vl_logic;
        HRDATA_RASBM_20 : out    vl_logic;
        HRDATA_RASBM_19 : out    vl_logic;
        HRDATA_RASBM_18 : out    vl_logic;
        HRDATA_RASBM_17 : out    vl_logic;
        HRDATA_RASBM_16 : out    vl_logic;
        HRDATA_RASBM_15 : out    vl_logic;
        HRDATA_RASBM_14 : out    vl_logic;
        HRDATA_RASBM_13 : out    vl_logic;
        HRDATA_RASBM_12 : out    vl_logic;
        HRDATA_RASBM_11 : out    vl_logic;
        HRDATA_RASBM_10 : out    vl_logic;
        HRDATA_RASBM_9  : out    vl_logic;
        HRDATA_RASBM_8  : out    vl_logic;
        HRDATA_RASBM_7  : out    vl_logic;
        HRDATA_RASBM_6  : out    vl_logic;
        HRDATA_RASBM_5  : out    vl_logic;
        HRDATA_RASBM_4  : out    vl_logic;
        HRDATA_RASBM_3  : out    vl_logic;
        HRDATA_RASBM_2  : out    vl_logic;
        HRDATA_RASBM_1  : out    vl_logic;
        HRDATA_RASBM_0  : out    vl_logic;
        HRESP_RASBM_1   : out    vl_logic;
        HRESP_RASBM_0   : out    vl_logic;
        HCLK_RASB       : out    vl_logic;
        HREADY_RASB     : out    vl_logic;
        HRESET_N_RASB   : out    vl_logic;
        RASB_DONE       : out    vl_logic;
        RASB_GSR_N      : out    vl_logic;
        RASB_IRQ_OUT    : out    vl_logic;
        EXT_CLK_P1_IN   : in     vl_logic;
        EXT_CLK_P2_IN   : in     vl_logic;
        EXT_DONE_IN     : in     vl_logic;
        QUAD_AND_FP0_7  : in     vl_logic;
        QUAD_AND_FP0_6  : in     vl_logic;
        QUAD_AND_FP0_5  : in     vl_logic;
        QUAD_AND_FP0_4  : in     vl_logic;
        QUAD_AND_FP0_3  : in     vl_logic;
        QUAD_AND_FP0_2  : in     vl_logic;
        QUAD_AND_FP0_1  : in     vl_logic;
        QUAD_AND_FP0_0  : in     vl_logic;
        QUAD_AND_FP1_7  : in     vl_logic;
        QUAD_AND_FP1_6  : in     vl_logic;
        QUAD_AND_FP1_5  : in     vl_logic;
        QUAD_AND_FP1_4  : in     vl_logic;
        QUAD_AND_FP1_3  : in     vl_logic;
        QUAD_AND_FP1_2  : in     vl_logic;
        QUAD_AND_FP1_1  : in     vl_logic;
        QUAD_AND_FP1_0  : in     vl_logic;
        QUAD_CLK_7      : in     vl_logic;
        QUAD_CLK_6      : in     vl_logic;
        QUAD_CLK_5      : in     vl_logic;
        QUAD_CLK_4      : in     vl_logic;
        QUAD_CLK_3      : in     vl_logic;
        QUAD_CLK_2      : in     vl_logic;
        QUAD_CLK_1      : in     vl_logic;
        QUAD_CLK_0      : in     vl_logic;
        QUAD_DONE_7     : in     vl_logic;
        QUAD_DONE_6     : in     vl_logic;
        QUAD_DONE_5     : in     vl_logic;
        QUAD_DONE_4     : in     vl_logic;
        QUAD_DONE_3     : in     vl_logic;
        QUAD_DONE_2     : in     vl_logic;
        QUAD_DONE_1     : in     vl_logic;
        QUAD_DONE_0     : in     vl_logic;
        QUAD_OR_FP0_7   : in     vl_logic;
        QUAD_OR_FP0_6   : in     vl_logic;
        QUAD_OR_FP0_5   : in     vl_logic;
        QUAD_OR_FP0_4   : in     vl_logic;
        QUAD_OR_FP0_3   : in     vl_logic;
        QUAD_OR_FP0_2   : in     vl_logic;
        QUAD_OR_FP0_1   : in     vl_logic;
        QUAD_OR_FP0_0   : in     vl_logic;
        QUAD_OR_FP1_7   : in     vl_logic;
        QUAD_OR_FP1_6   : in     vl_logic;
        QUAD_OR_FP1_5   : in     vl_logic;
        QUAD_OR_FP1_4   : in     vl_logic;
        QUAD_OR_FP1_3   : in     vl_logic;
        QUAD_OR_FP1_2   : in     vl_logic;
        QUAD_OR_FP1_1   : in     vl_logic;
        QUAD_OR_FP1_0   : in     vl_logic;
        QUAD_RST_N_7    : in     vl_logic;
        QUAD_RST_N_6    : in     vl_logic;
        QUAD_RST_N_5    : in     vl_logic;
        QUAD_RST_N_4    : in     vl_logic;
        QUAD_RST_N_3    : in     vl_logic;
        QUAD_RST_N_2    : in     vl_logic;
        QUAD_RST_N_1    : in     vl_logic;
        QUAD_RST_N_0    : in     vl_logic;
        QUAD_START_7    : in     vl_logic;
        QUAD_START_6    : in     vl_logic;
        QUAD_START_5    : in     vl_logic;
        QUAD_START_4    : in     vl_logic;
        QUAD_START_3    : in     vl_logic;
        QUAD_START_2    : in     vl_logic;
        QUAD_START_1    : in     vl_logic;
        QUAD_START_0    : in     vl_logic;
        EXT_CLK_P1_OUT  : out    vl_logic;
        EXT_CLK_P2_OUT  : out    vl_logic;
        EXT_DONE_OUT    : out    vl_logic;
        GRP_CLK_P1_L_3  : out    vl_logic;
        GRP_CLK_P1_L_2  : out    vl_logic;
        GRP_CLK_P1_L_1  : out    vl_logic;
        GRP_CLK_P1_L_0  : out    vl_logic;
        GRP_CLK_P2_L_3  : out    vl_logic;
        GRP_CLK_P2_L_2  : out    vl_logic;
        GRP_CLK_P2_L_1  : out    vl_logic;
        GRP_CLK_P2_L_0  : out    vl_logic;
        GRP_DESKEW_ERROR_L_3: out    vl_logic;
        GRP_DESKEW_ERROR_L_2: out    vl_logic;
        GRP_DESKEW_ERROR_L_1: out    vl_logic;
        GRP_DESKEW_ERROR_L_0: out    vl_logic;
        GRP_DONE_L_3    : out    vl_logic;
        GRP_DONE_L_2    : out    vl_logic;
        GRP_DONE_L_1    : out    vl_logic;
        GRP_DONE_L_0    : out    vl_logic;
        GRP_START_L_3   : out    vl_logic;
        GRP_START_L_2   : out    vl_logic;
        GRP_START_L_1   : out    vl_logic;
        GRP_START_L_0   : out    vl_logic;
        GRP_CLK_P1_R_3  : out    vl_logic;
        GRP_CLK_P1_R_2  : out    vl_logic;
        GRP_CLK_P1_R_1  : out    vl_logic;
        GRP_CLK_P1_R_0  : out    vl_logic;
        GRP_CLK_P2_R_3  : out    vl_logic;
        GRP_CLK_P2_R_2  : out    vl_logic;
        GRP_CLK_P2_R_1  : out    vl_logic;
        GRP_CLK_P2_R_0  : out    vl_logic;
        GRP_DESKEW_ERROR_R_3: out    vl_logic;
        GRP_DESKEW_ERROR_R_2: out    vl_logic;
        GRP_DESKEW_ERROR_R_1: out    vl_logic;
        GRP_DESKEW_ERROR_R_0: out    vl_logic;
        GRP_DONE_R_3    : out    vl_logic;
        GRP_DONE_R_2    : out    vl_logic;
        GRP_DONE_R_1    : out    vl_logic;
        GRP_DONE_R_0    : out    vl_logic;
        GRP_START_R_3   : out    vl_logic;
        GRP_START_R_2   : out    vl_logic;
        GRP_START_R_1   : out    vl_logic;
        GRP_START_R_0   : out    vl_logic;
        LPCS_INT_3      : in     vl_logic;
        LPCS_INT_2      : in     vl_logic;
        LPCS_INT_1      : in     vl_logic;
        LPCS_INT_0      : in     vl_logic;
        LPCS_RDATA_Q0_7 : in     vl_logic;
        LPCS_RDATA_Q0_6 : in     vl_logic;
        LPCS_RDATA_Q0_5 : in     vl_logic;
        LPCS_RDATA_Q0_4 : in     vl_logic;
        LPCS_RDATA_Q0_3 : in     vl_logic;
        LPCS_RDATA_Q0_2 : in     vl_logic;
        LPCS_RDATA_Q0_1 : in     vl_logic;
        LPCS_RDATA_Q0_0 : in     vl_logic;
        LPCS_RDATA_Q1_7 : in     vl_logic;
        LPCS_RDATA_Q1_6 : in     vl_logic;
        LPCS_RDATA_Q1_5 : in     vl_logic;
        LPCS_RDATA_Q1_4 : in     vl_logic;
        LPCS_RDATA_Q1_3 : in     vl_logic;
        LPCS_RDATA_Q1_2 : in     vl_logic;
        LPCS_RDATA_Q1_1 : in     vl_logic;
        LPCS_RDATA_Q1_0 : in     vl_logic;
        LPCS_RDATA_Q2_7 : in     vl_logic;
        LPCS_RDATA_Q2_6 : in     vl_logic;
        LPCS_RDATA_Q2_5 : in     vl_logic;
        LPCS_RDATA_Q2_4 : in     vl_logic;
        LPCS_RDATA_Q2_3 : in     vl_logic;
        LPCS_RDATA_Q2_2 : in     vl_logic;
        LPCS_RDATA_Q2_1 : in     vl_logic;
        LPCS_RDATA_Q2_0 : in     vl_logic;
        LPCS_RDATA_Q3_7 : in     vl_logic;
        LPCS_RDATA_Q3_6 : in     vl_logic;
        LPCS_RDATA_Q3_5 : in     vl_logic;
        LPCS_RDATA_Q3_4 : in     vl_logic;
        LPCS_RDATA_Q3_3 : in     vl_logic;
        LPCS_RDATA_Q3_2 : in     vl_logic;
        LPCS_RDATA_Q3_1 : in     vl_logic;
        LPCS_RDATA_Q3_0 : in     vl_logic;
        LPCS_ADDR_7     : out    vl_logic;
        LPCS_ADDR_6     : out    vl_logic;
        LPCS_ADDR_5     : out    vl_logic;
        LPCS_ADDR_4     : out    vl_logic;
        LPCS_ADDR_3     : out    vl_logic;
        LPCS_ADDR_2     : out    vl_logic;
        LPCS_ADDR_1     : out    vl_logic;
        LPCS_ADDR_0     : out    vl_logic;
        LPCS_WDATA_7    : out    vl_logic;
        LPCS_WDATA_6    : out    vl_logic;
        LPCS_WDATA_5    : out    vl_logic;
        LPCS_WDATA_4    : out    vl_logic;
        LPCS_WDATA_3    : out    vl_logic;
        LPCS_WDATA_2    : out    vl_logic;
        LPCS_WDATA_1    : out    vl_logic;
        LPCS_WDATA_0    : out    vl_logic;
        LPCS_C_15       : out    vl_logic;
        LPCS_C_14       : out    vl_logic;
        LPCS_C_13       : out    vl_logic;
        LPCS_C_12       : out    vl_logic;
        LPCS_C_11       : out    vl_logic;
        LPCS_C_10       : out    vl_logic;
        LPCS_C_9        : out    vl_logic;
        LPCS_C_8        : out    vl_logic;
        LPCS_C_7        : out    vl_logic;
        LPCS_C_6        : out    vl_logic;
        LPCS_C_5        : out    vl_logic;
        LPCS_C_4        : out    vl_logic;
        LPCS_C_3        : out    vl_logic;
        LPCS_C_2        : out    vl_logic;
        LPCS_C_1        : out    vl_logic;
        LPCS_C_0        : out    vl_logic;
        LPCS_Q_3        : out    vl_logic;
        LPCS_Q_2        : out    vl_logic;
        LPCS_Q_1        : out    vl_logic;
        LPCS_Q_0        : out    vl_logic;
        LPCS_RD         : out    vl_logic;
        LPCS_WSTB       : out    vl_logic;
        LPCS_QUAD_ID0_1 : out    vl_logic;
        LPCS_QUAD_ID0_0 : out    vl_logic;
        LPCS_QUAD_ID1_1 : out    vl_logic;
        LPCS_QUAD_ID1_0 : out    vl_logic;
        LPCS_QUAD_ID2_1 : out    vl_logic;
        LPCS_QUAD_ID2_0 : out    vl_logic;
        LPCS_QUAD_ID3_1 : out    vl_logic;
        LPCS_QUAD_ID3_0 : out    vl_logic;
        RPCS_INT_3      : in     vl_logic;
        RPCS_INT_2      : in     vl_logic;
        RPCS_INT_1      : in     vl_logic;
        RPCS_INT_0      : in     vl_logic;
        RPCS_RDATA_Q0_7 : in     vl_logic;
        RPCS_RDATA_Q0_6 : in     vl_logic;
        RPCS_RDATA_Q0_5 : in     vl_logic;
        RPCS_RDATA_Q0_4 : in     vl_logic;
        RPCS_RDATA_Q0_3 : in     vl_logic;
        RPCS_RDATA_Q0_2 : in     vl_logic;
        RPCS_RDATA_Q0_1 : in     vl_logic;
        RPCS_RDATA_Q0_0 : in     vl_logic;
        RPCS_RDATA_Q1_7 : in     vl_logic;
        RPCS_RDATA_Q1_6 : in     vl_logic;
        RPCS_RDATA_Q1_5 : in     vl_logic;
        RPCS_RDATA_Q1_4 : in     vl_logic;
        RPCS_RDATA_Q1_3 : in     vl_logic;
        RPCS_RDATA_Q1_2 : in     vl_logic;
        RPCS_RDATA_Q1_1 : in     vl_logic;
        RPCS_RDATA_Q1_0 : in     vl_logic;
        RPCS_RDATA_Q2_7 : in     vl_logic;
        RPCS_RDATA_Q2_6 : in     vl_logic;
        RPCS_RDATA_Q2_5 : in     vl_logic;
        RPCS_RDATA_Q2_4 : in     vl_logic;
        RPCS_RDATA_Q2_3 : in     vl_logic;
        RPCS_RDATA_Q2_2 : in     vl_logic;
        RPCS_RDATA_Q2_1 : in     vl_logic;
        RPCS_RDATA_Q2_0 : in     vl_logic;
        RPCS_RDATA_Q3_7 : in     vl_logic;
        RPCS_RDATA_Q3_6 : in     vl_logic;
        RPCS_RDATA_Q3_5 : in     vl_logic;
        RPCS_RDATA_Q3_4 : in     vl_logic;
        RPCS_RDATA_Q3_3 : in     vl_logic;
        RPCS_RDATA_Q3_2 : in     vl_logic;
        RPCS_RDATA_Q3_1 : in     vl_logic;
        RPCS_RDATA_Q3_0 : in     vl_logic;
        RPCS_ADDR_7     : out    vl_logic;
        RPCS_ADDR_6     : out    vl_logic;
        RPCS_ADDR_5     : out    vl_logic;
        RPCS_ADDR_4     : out    vl_logic;
        RPCS_ADDR_3     : out    vl_logic;
        RPCS_ADDR_2     : out    vl_logic;
        RPCS_ADDR_1     : out    vl_logic;
        RPCS_ADDR_0     : out    vl_logic;
        RPCS_WDATA_7    : out    vl_logic;
        RPCS_WDATA_6    : out    vl_logic;
        RPCS_WDATA_5    : out    vl_logic;
        RPCS_WDATA_4    : out    vl_logic;
        RPCS_WDATA_3    : out    vl_logic;
        RPCS_WDATA_2    : out    vl_logic;
        RPCS_WDATA_1    : out    vl_logic;
        RPCS_WDATA_0    : out    vl_logic;
        RPCS_C_15       : out    vl_logic;
        RPCS_C_14       : out    vl_logic;
        RPCS_C_13       : out    vl_logic;
        RPCS_C_12       : out    vl_logic;
        RPCS_C_11       : out    vl_logic;
        RPCS_C_10       : out    vl_logic;
        RPCS_C_9        : out    vl_logic;
        RPCS_C_8        : out    vl_logic;
        RPCS_C_7        : out    vl_logic;
        RPCS_C_6        : out    vl_logic;
        RPCS_C_5        : out    vl_logic;
        RPCS_C_4        : out    vl_logic;
        RPCS_C_3        : out    vl_logic;
        RPCS_C_2        : out    vl_logic;
        RPCS_C_1        : out    vl_logic;
        RPCS_C_0        : out    vl_logic;
        RPCS_Q_3        : out    vl_logic;
        RPCS_Q_2        : out    vl_logic;
        RPCS_Q_1        : out    vl_logic;
        RPCS_Q_0        : out    vl_logic;
        RPCS_RD         : out    vl_logic;
        RPCS_WSTB       : out    vl_logic;
        RPCS_QUAD_ID0_1 : out    vl_logic;
        RPCS_QUAD_ID0_0 : out    vl_logic;
        RPCS_QUAD_ID1_1 : out    vl_logic;
        RPCS_QUAD_ID1_0 : out    vl_logic;
        RPCS_QUAD_ID2_1 : out    vl_logic;
        RPCS_QUAD_ID2_0 : out    vl_logic;
        RPCS_QUAD_ID3_1 : out    vl_logic;
        RPCS_QUAD_ID3_0 : out    vl_logic;
        DMA_RD_DATA_31  : in     vl_logic;
        DMA_RD_DATA_30  : in     vl_logic;
        DMA_RD_DATA_29  : in     vl_logic;
        DMA_RD_DATA_28  : in     vl_logic;
        DMA_RD_DATA_27  : in     vl_logic;
        DMA_RD_DATA_26  : in     vl_logic;
        DMA_RD_DATA_25  : in     vl_logic;
        DMA_RD_DATA_24  : in     vl_logic;
        DMA_RD_DATA_23  : in     vl_logic;
        DMA_RD_DATA_22  : in     vl_logic;
        DMA_RD_DATA_21  : in     vl_logic;
        DMA_RD_DATA_20  : in     vl_logic;
        DMA_RD_DATA_19  : in     vl_logic;
        DMA_RD_DATA_18  : in     vl_logic;
        DMA_RD_DATA_17  : in     vl_logic;
        DMA_RD_DATA_16  : in     vl_logic;
        DMA_RD_DATA_15  : in     vl_logic;
        DMA_RD_DATA_14  : in     vl_logic;
        DMA_RD_DATA_13  : in     vl_logic;
        DMA_RD_DATA_12  : in     vl_logic;
        DMA_RD_DATA_11  : in     vl_logic;
        DMA_RD_DATA_10  : in     vl_logic;
        DMA_RD_DATA_9   : in     vl_logic;
        DMA_RD_DATA_8   : in     vl_logic;
        DMA_RD_DATA_7   : in     vl_logic;
        DMA_RD_DATA_6   : in     vl_logic;
        DMA_RD_DATA_5   : in     vl_logic;
        DMA_RD_DATA_4   : in     vl_logic;
        DMA_RD_DATA_3   : in     vl_logic;
        DMA_RD_DATA_2   : in     vl_logic;
        DMA_RD_DATA_1   : in     vl_logic;
        DMA_RD_DATA_0   : in     vl_logic;
        DMA_RD_PARITY_3 : in     vl_logic;
        DMA_RD_PARITY_2 : in     vl_logic;
        DMA_RD_PARITY_1 : in     vl_logic;
        DMA_RD_PARITY_0 : in     vl_logic;
        DMA_RETRY       : in     vl_logic;
        DMA_TA          : in     vl_logic;
        DMA_TEA         : in     vl_logic;
        DMA_TRI_CTL     : in     vl_logic;
        DMA_TRI_DATA    : in     vl_logic
    );
end SYSBUSA_sim;
