library verilog;
use verilog.vl_types.all;
entity pcs_quad_clocks is
    port(
        txclk0          : in     vl_logic;
        txclk1          : in     vl_logic;
        txclk2          : in     vl_logic;
        txclk3          : in     vl_logic;
        test_clk        : in     vl_logic;
        lane_tx_rst0    : in     vl_logic;
        lane_tx_rst1    : in     vl_logic;
        lane_tx_rst2    : in     vl_logic;
        lane_tx_rst3    : in     vl_logic;
        lane_rx_rst0    : in     vl_logic;
        lane_rx_rst1    : in     vl_logic;
        lane_rx_rst2    : in     vl_logic;
        lane_rx_rst3    : in     vl_logic;
        ffc_lane_tx_rst0: in     vl_logic;
        ffc_lane_tx_rst1: in     vl_logic;
        ffc_lane_tx_rst2: in     vl_logic;
        ffc_lane_tx_rst3: in     vl_logic;
        ffc_lane_rx_rst0: in     vl_logic;
        ffc_lane_rx_rst1: in     vl_logic;
        ffc_lane_rx_rst2: in     vl_logic;
        ffc_lane_rx_rst3: in     vl_logic;
        ffc_quad_rst    : in     vl_logic;
        ffc_macro_rst   : in     vl_logic;
        pwrupres        : in     vl_logic;
        qif_quad_rst    : in     vl_logic;
        qif_macro_rst   : in     vl_logic;
        fpga_reset_en   : in     vl_logic;
        rxclk0          : in     vl_logic;
        rxclk1          : in     vl_logic;
        rxclk2          : in     vl_logic;
        rxclk3          : in     vl_logic;
        cascade_clk     : in     vl_logic;
        sysclk0         : out    vl_logic;
        sysclk1         : out    vl_logic;
        sysclk2         : out    vl_logic;
        sysclk3         : out    vl_logic;
        sys_txrst0_n    : out    vl_logic;
        sys_txrst1_n    : out    vl_logic;
        sys_txrst2_n    : out    vl_logic;
        sys_txrst3_n    : out    vl_logic;
        sys_rxrst0_n    : out    vl_logic;
        sys_rxrst1_n    : out    vl_logic;
        sys_rxrst2_n    : out    vl_logic;
        sys_rxrst3_n    : out    vl_logic;
        pcs_rxclk0      : out    vl_logic;
        pcs_rxrst0_n    : out    vl_logic;
        pcs_rxclk1      : out    vl_logic;
        pcs_rxrst1_n    : out    vl_logic;
        pcs_rxclk2      : out    vl_logic;
        pcs_rxrst2_n    : out    vl_logic;
        pcs_rxclk3      : out    vl_logic;
        pcs_rxrst3_n    : out    vl_logic;
        m_rxclk0        : out    vl_logic;
        m_rxrst0_n      : out    vl_logic;
        m_rxclk1        : out    vl_logic;
        m_rxrst1_n      : out    vl_logic;
        m_rxclk2        : out    vl_logic;
        m_rxrst2_n      : out    vl_logic;
        m_rxclk3        : out    vl_logic;
        m_rxrst3_n      : out    vl_logic;
        fb_rxclk0       : out    vl_logic;
        fb_rxrst0_n     : out    vl_logic;
        fb_rxclk1       : out    vl_logic;
        fb_rxrst1_n     : out    vl_logic;
        fb_rxclk2       : out    vl_logic;
        fb_rxrst2_n     : out    vl_logic;
        fb_rxclk3       : out    vl_logic;
        fb_rxrst3_n     : out    vl_logic;
        ff_sysclk_p1    : out    vl_logic;
        ff_sysclk0      : out    vl_logic;
        ff_sysclk1      : out    vl_logic;
        ff_sysclk2      : out    vl_logic;
        ff_sysclk3      : out    vl_logic;
        ff_rxclk_p1     : out    vl_logic;
        ff_rxclk_p2     : out    vl_logic;
        ff_rxclk0       : out    vl_logic;
        ff_rxclk1       : out    vl_logic;
        ff_rxclk2       : out    vl_logic;
        ff_rxclk3       : out    vl_logic;
        quad_clk        : out    vl_logic;
        pwr_on_rst      : out    vl_logic;
        macrorst        : out    vl_logic;
        rst_n           : out    vl_logic;
        scan_mode       : in     vl_logic;
        scan_rstn       : in     vl_logic;
        test_mode       : in     vl_logic_vector(2 downto 0);
        fb_tx_mode      : in     vl_logic;
        fb_rx_mode      : in     vl_logic;
        uc_mode         : in     vl_logic;
        pcs_mode        : in     vl_logic;
        x4_mode         : in     vl_logic;
        cascade_en      : in     vl_logic;
        mclksel_0       : in     vl_logic_vector(1 downto 0);
        mclksel_1       : in     vl_logic_vector(1 downto 0);
        mclksel_2       : in     vl_logic_vector(1 downto 0);
        mclksel_3       : in     vl_logic_vector(1 downto 0);
        qclksel         : in     vl_logic_vector(1 downto 0);
        ff_sysclk_p1_sel: in     vl_logic_vector(1 downto 0);
        ff_rxclk_p1_sel : in     vl_logic_vector(1 downto 0);
        ff_rxclk_p2_sel : in     vl_logic_vector(1 downto 0);
        sb_loopback_0   : in     vl_logic;
        sb_loopback_1   : in     vl_logic;
        sb_loopback_2   : in     vl_logic;
        sb_loopback_3   : in     vl_logic;
        TIE_HIGH        : out    vl_logic;
        TIE_LOW         : out    vl_logic
    );
end pcs_quad_clocks;
