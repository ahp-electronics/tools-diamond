library verilog;
use verilog.vl_types.all;
entity e2_serdes_ch_model is
    port(
        HDINPi          : in     vl_logic;
        HDINNi          : in     vl_logic;
        ck_core_rx      : in     vl_logic;
        rx_refck_local  : in     vl_logic;
        ck3g4tx         : in     vl_logic;
        mrstb           : in     vl_logic;
        rpwdnb          : in     vl_logic;
        tpwdnb          : in     vl_logic;
        rrst            : in     vl_logic;
        tdi             : in     vl_logic_vector(9 downto 0);
        oob_en          : in     vl_logic;
        pci_en          : in     vl_logic;
        pci_ei_en       : in     vl_logic;
        pci_det_en      : in     vl_logic;
        pci_det_ct      : in     vl_logic;
        bs2pad          : in     vl_logic;
        bstxsel         : in     vl_logic;
        bsrxsel         : in     vl_logic;
        auto_calib_enb  : in     vl_logic;
        auto_facq_enb   : in     vl_logic;
        band_threshold  : in     vl_logic_vector(5 downto 0);
        bus8bit_sel     : in     vl_logic;
        calib_ck_mode   : in     vl_logic;
        calib_time_sel  : in     vl_logic_vector(1 downto 0);
        cdr_lol_set     : in     vl_logic_vector(1 downto 0);
        dac_bdavoid_enb : in     vl_logic;
        fc2dco_dloop    : in     vl_logic;
        lb_ctl          : in     vl_logic_vector(3 downto 0);
        pd_i_set        : in     vl_logic_vector(1 downto 0);
        rate_mode_rx    : in     vl_logic;
        rate_mode_tx    : in     vl_logic;
        rcv_dcc_en      : in     vl_logic;
        refck25x        : in     vl_logic;
        refck_mode      : in     vl_logic_vector(1 downto 0);
        reg_band_offset : in     vl_logic_vector(3 downto 0);
        reg_band_range  : in     vl_logic_vector(2 downto 0);
        reg_band_sel    : in     vl_logic_vector(5 downto 0);
        reg_calib_rst   : in     vl_logic;
        reg_facq_rst    : in     vl_logic;
        reg_idac_en     : in     vl_logic;
        reg_idac_sel    : in     vl_logic_vector(9 downto 0);
        req_en          : in     vl_logic;
        req_i_set       : in     vl_logic_vector(2 downto 0);
        req_lvl_set     : in     vl_logic;
        rlos_hset       : in     vl_logic_vector(2 downto 0);
        rlos_lset       : in     vl_logic_vector(2 downto 0);
        rterm_rx        : in     vl_logic_vector(1 downto 0);
        rterm_rxadj     : in     vl_logic_vector(1 downto 0);
        rterm_tx        : in     vl_logic_vector(1 downto 0);
        rx_dco_ck_div   : in     vl_logic_vector(2 downto 0);
        rx_refck_sel    : in     vl_logic_vector(1 downto 0);
        tdrv_amp        : in     vl_logic_vector(2 downto 0);
        tdrv_dat_sel    : in     vl_logic_vector(1 downto 0);
        tdrv_pre_en     : in     vl_logic;
        tdrv_pre_set    : in     vl_logic_vector(2 downto 0);
        HDOUTPi         : out    vl_logic;
        HDOUTNi         : out    vl_logic;
        pci_connect     : out    vl_logic;
        pci_det_done    : out    vl_logic;
        rdi             : out    vl_logic_vector(9 downto 0);
        rcki            : out    vl_logic;
        rlol            : out    vl_logic;
        rlos_lo         : out    vl_logic;
        rlos_hi         : out    vl_logic;
        tcki            : out    vl_logic;
        dco_calib_done  : out    vl_logic;
        dco_calib_err   : out    vl_logic;
        dco_facq_done   : out    vl_logic;
        dco_facq_err    : out    vl_logic;
        dco_status      : out    vl_logic_vector(15 downto 0);
        oob_out         : out    vl_logic;
        bs4pad          : out    vl_logic
    );
end e2_serdes_ch_model;
