library verilog;
use verilog.vl_types.all;
entity delc0p5x2v1mce is
    port(
        A               : in     vl_logic;
        Z               : out    vl_logic
    );
end delc0p5x2v1mce;
