library verilog;
use verilog.vl_types.all;
entity sys_bus_top is
    generic(
        QUAD            : integer := 8;
        GRP             : integer := 4
    );
    port(
        USER_IRQ_OUT    : out    vl_logic;
        UPDTDR_RASB     : out    vl_logic;
        UPDTDR_LASB     : out    vl_logic;
        UPDTBSR         : out    vl_logic;
        TRI_ION         : out    vl_logic;
        TRESET_RASB     : out    vl_logic;
        TRESET_LASB     : out    vl_logic;
        TRESET          : out    vl_logic;
        TMS_CIB         : out    vl_logic;
        TDOEN           : out    vl_logic;
        TDOE            : out    vl_logic;
        TDO             : out    vl_logic;
        TDI_CIB         : out    vl_logic;
        TDI1_RASB       : out    vl_logic;
        TDI1_LASB       : out    vl_logic;
        TCK_CIB         : out    vl_logic;
        TCK2_RASB       : out    vl_logic;
        TCK2_LASB       : out    vl_logic;
        TCK2            : out    vl_logic;
        SYSB_DEBUG      : out    vl_logic_vector(23 downto 0);
        SRI_WR          : out    vl_logic;
        SRI_WDATA       : out    vl_logic;
        SRI_RST_N       : out    vl_logic;
        SRI_RD          : out    vl_logic;
        SRI_CLK         : out    vl_logic;
        SRI_ADDR        : out    vl_logic_vector(9 downto 0);
        SPI_TRI_ION     : out    vl_logic;
        SHIFT_ADDR_2ND  : out    vl_logic;
        SHIFT_ADDR_1ST  : out    vl_logic;
        SHDR_RASB       : out    vl_logic;
        SHDR_LASB       : out    vl_logic;
        SHBSRN          : out    vl_logic;
        SERIAL_DATA     : out    vl_logic;
        SCANEN_RASB     : out    vl_logic;
        SCANEN_LASB     : out    vl_logic;
        SBWR_O          : out    vl_logic_vector(33 downto 0);
        RUNTST_RASB     : out    vl_logic;
        RUNTST_LASB     : out    vl_logic;
        RST_DATA_REG_N  : out    vl_logic;
        RST_ADDR_REG    : out    vl_logic;
        RPCS_WSTB       : out    vl_logic;
        RPCS_Q          : out    vl_logic_vector(3 downto 0);
        RPCS_C          : out    vl_logic_vector(15 downto 0);
        RDY_BUSY_N      : out    vl_logic;
        RDBK_DATA       : out    vl_logic;
        RASB_PWRUPRES   : out    vl_logic;
        RASB_IRQ_OUT    : out    vl_logic;
        RASB_GSR_N      : out    vl_logic;
        RASB_DONE       : out    vl_logic;
        QOUT            : out    vl_logic;
        Q15_LOCAL_RDATA : out    vl_logic_vector(7 downto 0);
        PWR_ON          : out    vl_logic;
        PWRUPRES        : out    vl_logic;
        PSRTRST         : out    vl_logic;
        PSRSFTN         : out    vl_logic;
        PSRENABLE3      : out    vl_logic;
        PSRENABLE2      : out    vl_logic;
        PSRENABLE1      : out    vl_logic;
        PSRCAP          : out    vl_logic;
        PRDY_TS         : out    vl_logic;
        PD7_3_TS        : out    vl_logic;
        PD31_16_TS      : out    vl_logic;
        PD2_0_TS        : out    vl_logic;
        PD15_8_TS       : out    vl_logic;
        PCS_TRI_ION     : out    vl_logic;
        PCS_M_TRI_ION   : out    vl_logic;
        PA_OUT          : out    vl_logic_vector(21 downto 0);
        PAD_DONE        : out    vl_logic;
        MPI_TRI_ION     : out    vl_logic_vector(2 downto 0);
        MPI_IRQ_N       : out    vl_logic;
        MPI_DP_TS       : out    vl_logic_vector(2 downto 0);
        MPI_DP_TRI_ION  : out    vl_logic_vector(2 downto 0);
        MPI_CNTL_TS     : out    vl_logic;
        MPC_TEA         : out    vl_logic;
        MPC_TA          : out    vl_logic;
        MPC_RETRY       : out    vl_logic;
        MPC_RD_PARITY   : out    vl_logic_vector(0 to 3);
        MPC_RD_DATA     : out    vl_logic_vector(0 to 31);
        LPCS_WSTB       : out    vl_logic;
        LPCS_WDATA      : out    vl_logic_vector(7 downto 0);
        LPCS_RD         : out    vl_logic;
        LPCS_Q          : out    vl_logic_vector(3 downto 0);
        LPCS_C          : out    vl_logic_vector(15 downto 0);
        LPCS_ADDR       : out    vl_logic_vector(7 downto 0);
        LD_RDBKD        : out    vl_logic;
        LDC_N           : out    vl_logic;
        LASB_PWRUPRES   : out    vl_logic;
        LASB_IRQ_OUT    : out    vl_logic;
        LASB_GSR_N      : out    vl_logic;
        LASB_DONE       : out    vl_logic;
        JUPDATE         : out    vl_logic;
        JTDI            : out    vl_logic;
        JTCK            : out    vl_logic;
        JSHIFT          : out    vl_logic;
        JSCANIN         : out    vl_logic;
        JSCANENABLE     : out    vl_logic_vector(8 downto 1);
        JRTI            : out    vl_logic_vector(8 downto 1);
        JRSTN           : out    vl_logic;
        JCE             : out    vl_logic_vector(8 downto 1);
        IS_SLAVE3_OUT   : out    vl_logic;
        IS_SLAVE2_OUT   : out    vl_logic;
        IS_SLAVE1_OUT   : out    vl_logic;
        IS_SLAVE0_OUT   : out    vl_logic;
        IQA_TX_ALIGN_R  : out    vl_logic;
        IQA_TX_ALIGN_L  : out    vl_logic;
        INTEST          : out    vl_logic;
        INIT_N          : out    vl_logic;
        INIT_1_DATA     : out    vl_logic;
        HRESP_RASBM     : out    vl_logic_vector(1 downto 0);
        HRESP_LASBM     : out    vl_logic_vector(1 downto 0);
        HRESET_N_RASB   : out    vl_logic;
        HRESET_N_LASB   : out    vl_logic;
        HREADY_RASB     : out    vl_logic;
        HREADY_LASB     : out    vl_logic;
        HRDATA_RASBM    : out    vl_logic_vector(35 downto 0);
        HRDATA_LASBM    : out    vl_logic_vector(35 downto 0);
        HIGHZ           : out    vl_logic;
        HGRANT_RASBM    : out    vl_logic;
        HGRANT_LASBM    : out    vl_logic;
        HDC             : out    vl_logic;
        HCLK_CIB        : out    vl_logic;
        GSR_N           : out    vl_logic;
        GSRN_SYNC       : out    vl_logic;
        GRP3_WRST_OUT_N : out    vl_logic;
        GRP3_RRST_OUT_N : out    vl_logic;
        GRP2_WRST_OUT_N : out    vl_logic;
        GRP2_RRST_OUT_N : out    vl_logic;
        GRP1_WRST_OUT_N : out    vl_logic;
        GRP1_RRST_OUT_N : out    vl_logic;
        GRP0_WRST_OUT_N : out    vl_logic;
        GRP0_RRST_OUT_N : out    vl_logic;
        GOT_DATA        : out    vl_logic;
        GOT_ADDR        : out    vl_logic;
        FSWRN           : out    vl_logic;
        FSWDATA         : out    vl_logic_vector(35 downto 0);
        FSSIZE          : out    vl_logic_vector(1 downto 0);
        FSRDY           : out    vl_logic;
        FSADDR          : out    vl_logic_vector(17 downto 0);
        FMRETRY         : out    vl_logic;
        FMRDATA         : out    vl_logic_vector(35 downto 0);
        FMERR           : out    vl_logic;
        FMACK           : out    vl_logic;
        EXT_DONE_OUT    : out    vl_logic;
        EXT_CLK_P2_OUT  : out    vl_logic;
        EXT_CLK_P1_OUT  : out    vl_logic;
        EN_OSC          : out    vl_logic;
        EN_CCLK_N       : out    vl_logic;
        EN_ADDR_INCR    : out    vl_logic;
        EN_ADDR         : out    vl_logic;
        DOUT            : out    vl_logic;
        DONE            : out    vl_logic;
        DOBIST_RASB     : out    vl_logic;
        DOBIST_LASB     : out    vl_logic;
        DEBUG_BUS       : out    vl_logic_vector(15 downto 0);
        CPTDR_RASB      : out    vl_logic;
        CPTDR_LASB      : out    vl_logic;
        CPTBSR          : out    vl_logic;
        CFG_DATA_WR     : out    vl_logic;
        CFG_DATA_PC     : out    vl_logic;
        CFG_DATA        : out    vl_logic_vector(7 downto 0);
        CFG_CK          : out    vl_logic;
        CCLK_OUT        : out    vl_logic;
        CCLK_AD         : out    vl_logic;
        BS_MODE         : out    vl_logic;
        ADDR_TS         : out    vl_logic;
        GRP_CLK_P1_L    : out    vl_logic_vector;
        GRP_CLK_P2_L    : out    vl_logic_vector;
        GRP_DESKEW_ERROR_L: out    vl_logic_vector;
        GRP_DONE_L      : out    vl_logic_vector;
        GRP_START_L     : out    vl_logic_vector;
        GRP_CLK_P1_R    : out    vl_logic_vector;
        GRP_CLK_P2_R    : out    vl_logic_vector;
        GRP_DESKEW_ERROR_R: out    vl_logic_vector;
        GRP_DONE_R      : out    vl_logic_vector;
        GRP_START_R     : out    vl_logic_vector;
        HCLK_LASB       : out    vl_logic;
        HCLK_RASB       : out    vl_logic;
        RPCS_ADDR       : out    vl_logic_vector(7 downto 0);
        RPCS_RD         : out    vl_logic;
        RPCS_WDATA      : out    vl_logic_vector(7 downto 0);
        SYS_TRI_ION     : out    vl_logic;
        SYS_LOW         : out    vl_logic;
        SYS_HIGH        : out    vl_logic;
        PCS_LOW         : out    vl_logic;
        PCS_HIGH        : out    vl_logic;
        TDI1            : out    vl_logic;
        EN_PDWN         : out    vl_logic;
        WR_N            : in     vl_logic;
        USR_TDO         : in     vl_logic;
        USR_START_CLK   : in     vl_logic;
        USR_GSR         : in     vl_logic;
        USR_CLK         : in     vl_logic;
        USER_IRQ_IN     : in     vl_logic;
        TX_ALIGN        : in     vl_logic;
        TS_ALL          : in     vl_logic;
        TMS             : in     vl_logic;
        TDI             : in     vl_logic;
        TCK             : in     vl_logic;
        SYS_SE          : in     vl_logic;
        SYS_RST_N       : in     vl_logic;
        SRI_RDATA       : in     vl_logic_vector(63 downto 0);
        SO_BIST_RASB    : in     vl_logic;
        SO_BIST_LASB    : in     vl_logic;
        SED_CLK         : in     vl_logic;
        SCANOUT_RASB    : in     vl_logic;
        SCANOUT_LASB    : in     vl_logic;
        RPCS_RDATA      : in     vl_logic_vector(7 downto 0);
        RD_N            : in     vl_logic;
        RD_CFG_USR      : in     vl_logic;
        RD_CFG          : in     vl_logic;
        RDBK_ZERO_ALL_N : in     vl_logic;
        RDBK_DOUT       : in     vl_logic_vector(7 downto 0);
        RASB_SLAVE_ENABLE: in     vl_logic;
        RASB_SEL        : in     vl_logic;
        RASB_IRQ_MASTER : in     vl_logic;
        RASB_GSR        : in     vl_logic;
        RASB_CLK        : in     vl_logic;
        QUAD_START      : in     vl_logic_vector;
        QUAD_RST_N      : in     vl_logic_vector;
        QUAD_OR_FP1     : in     vl_logic_vector;
        QUAD_OR_FP0     : in     vl_logic_vector;
        QUAD_DONE       : in     vl_logic_vector;
        QUAD_CLK        : in     vl_logic_vector;
        QUAD_AND_FP1    : in     vl_logic_vector;
        QUAD_AND_FP0    : in     vl_logic_vector;
        PWRUP_NPUR      : in     vl_logic;
        PWRUP_E9        : in     vl_logic;
        PTEST_N         : in     vl_logic;
        PSROUT3         : in     vl_logic;
        PSROUT2         : in     vl_logic;
        PSROUT1         : in     vl_logic;
        PARTID          : in     vl_logic_vector(31 downto 0);
        MPI_RST_N       : in     vl_logic;
        MPI_CLK         : in     vl_logic;
        MPC_WR_PARITY   : in     vl_logic_vector(0 to 3);
        MPC_WR_DATA     : in     vl_logic_vector(0 to 31);
        MPC_TSIZ        : in     vl_logic_vector(0 to 1);
        MPC_BURST       : in     vl_logic;
        MPC_BDIP        : in     vl_logic;
        MPC_ADDR        : in     vl_logic_vector(14 to 31);
        MODE            : in     vl_logic_vector(3 downto 0);
        MC1_USR_TDO     : in     vl_logic;
        MC1_USR_SL      : in     vl_logic_vector(1 downto 0);
        MC1_USR_MR      : in     vl_logic_vector(1 downto 0);
        MC1_USR_CLK     : in     vl_logic;
        MC1_USERBIT     : in     vl_logic_vector(31 downto 0);
        MC1_USER        : in     vl_logic;
        MC1_TRI         : in     vl_logic_vector(3 downto 0);
        MC1_TIMEOUT_INDEX2: in     vl_logic_vector(3 downto 0);
        MC1_TIMEOUT_INDEX1: in     vl_logic_vector(3 downto 0);
        MC1_TEST_CTR    : in     vl_logic;
        MC1_SYS_RST     : in     vl_logic;
        MC1_STRT        : in     vl_logic_vector(4 downto 0);
        MC1_SPI_ADDR    : in     vl_logic_vector(31 downto 0);
        MC1_SED_CLK     : in     vl_logic;
        MC1_SCLK        : in     vl_logic;
        MC1_SCAN        : in     vl_logic_vector(8 downto 1);
        MC1_RST_RAM_N   : in     vl_logic;
        MC1_RST_HCLK_N  : in     vl_logic;
        MC1_RST_GSRN    : in     vl_logic;
        MC1_RST_BUS_N   : in     vl_logic;
        MC1_RDBK_REG    : in     vl_logic;
        MC1_PRIORITY_MPI: in     vl_logic_vector(1 downto 0);
        MC1_PRIORITY_FPGA: in     vl_logic_vector(1 downto 0);
        MC1_PRIORITY_ASB: in     vl_logic_vector(1 downto 0);
        MC1_PAR_ODD     : in     vl_logic;
        MC1_OSC_DIV     : in     vl_logic_vector(2 downto 0);
        MC1_OSC_CLK     : in     vl_logic;
        MC1_MPI_RST     : in     vl_logic;
        MC1_MPI_CLK     : in     vl_logic;
        MC1_MPI_ASYNC   : in     vl_logic;
        MC1_MPI         : in     vl_logic;
        MC1_MODE        : in     vl_logic_vector(3 downto 0);
        MC1_INTERRUPT_VECTOR_6: in     vl_logic_vector(31 downto 0);
        MC1_INTERRUPT_VECTOR_5: in     vl_logic_vector(31 downto 0);
        MC1_INTERRUPT_VECTOR_4: in     vl_logic_vector(31 downto 0);
        MC1_INTERRUPT_VECTOR_3: in     vl_logic_vector(31 downto 0);
        MC1_INTERRUPT_VECTOR_2: in     vl_logic_vector(31 downto 0);
        MC1_INTERRUPT_VECTOR_1: in     vl_logic_vector(31 downto 0);
        MC1_GSRN_SYNC   : in     vl_logic;
        MC1_GSRN_INV    : in     vl_logic;
        MC1_FPSC_CLK    : in     vl_logic;
        MC1_FPSC        : in     vl_logic;
        MC1_EXT_CCLK    : in     vl_logic;
        MC1_EN_SPI_N    : in     vl_logic;
        MC1_EN_SED      : in     vl_logic;
        MC1_EN_RDBK     : in     vl_logic;
        MC1_EN_OSC      : in     vl_logic;
        MC1_EN_ONCE     : in     vl_logic;
        MC1_EN_MPI_PARITY: in     vl_logic;
        MC1_DONE        : in     vl_logic_vector(1 downto 0);
        MC1_DIS_MODES   : in     vl_logic;
        LPCS_RDATA      : in     vl_logic_vector(7 downto 0);
        LAST_ADDR       : in     vl_logic_vector(13 downto 0);
        LASB_SLAVE_ENABLE: in     vl_logic;
        LASB_IRQ_MASTER : in     vl_logic;
        LASB_GSR        : in     vl_logic;
        LASB_CLK        : in     vl_logic;
        JTDO            : in     vl_logic_vector(8 downto 1);
        IS_SLAVE3_IN    : in     vl_logic;
        IS_SLAVE2_IN    : in     vl_logic;
        IS_SLAVE1_IN    : in     vl_logic;
        IS_SLAVE0_IN    : in     vl_logic;
        INITIN_N        : in     vl_logic;
        HWRITE_RASBM    : in     vl_logic;
        HWRITE_LASBM    : in     vl_logic;
        HWDATA_RASBM    : in     vl_logic_vector(35 downto 0);
        HWDATA_LASBM    : in     vl_logic_vector(35 downto 0);
        HTRANS_RASBM    : in     vl_logic_vector(1 downto 0);
        HTRANS_LASBM    : in     vl_logic_vector(1 downto 0);
        HSIZE_RASBM     : in     vl_logic_vector(1 downto 0);
        HSIZE_LASBM     : in     vl_logic_vector(1 downto 0);
        HLOCK_RASBM     : in     vl_logic;
        HLOCK_LASBM     : in     vl_logic;
        HBUSREQ_RASBM   : in     vl_logic;
        HBUSREQ_LASBM   : in     vl_logic;
        HBURST_RASBM    : in     vl_logic;
        HBURST_LASBM    : in     vl_logic;
        HADDR_RASBM     : in     vl_logic_vector(17 downto 0);
        HADDR_LASBM     : in     vl_logic_vector(17 downto 0);
        GRP3_WRST_IN_N  : in     vl_logic;
        GRP3_RRST_IN_N  : in     vl_logic;
        GRP2_WRST_IN_N  : in     vl_logic;
        GRP2_RRST_IN_N  : in     vl_logic;
        GRP1_WRST_IN_N  : in     vl_logic;
        GRP1_RRST_IN_N  : in     vl_logic;
        GRP0_WRST_IN_N  : in     vl_logic;
        GRP0_RRST_IN_N  : in     vl_logic;
        FSRETRY         : in     vl_logic;
        FSRESET_N       : in     vl_logic;
        FSRDATA         : in     vl_logic_vector(35 downto 0);
        FSIRQ           : in     vl_logic;
        FSERR           : in     vl_logic;
        FSCLK           : in     vl_logic;
        FSACK           : in     vl_logic;
        FMWRN           : in     vl_logic;
        FMWDATA         : in     vl_logic_vector(35 downto 0);
        FMSIZE          : in     vl_logic_vector(1 downto 0);
        FMRESET_N       : in     vl_logic;
        FMRDY           : in     vl_logic;
        FMLOCK          : in     vl_logic;
        FMIRQ           : in     vl_logic;
        FMCLK           : in     vl_logic;
        FMBURST         : in     vl_logic;
        FMADDR          : in     vl_logic_vector(17 downto 0);
        EXT_DONE_IN     : in     vl_logic;
        EXT_CLK_P2_IN   : in     vl_logic;
        EXT_CLK_P1_IN   : in     vl_logic;
        DONEIN          : in     vl_logic;
        DMA_TRI_DATA    : in     vl_logic;
        DMA_TRI_CTL     : in     vl_logic;
        DMA_TEA         : in     vl_logic;
        DMA_TA          : in     vl_logic;
        DMA_RETRY       : in     vl_logic;
        DMA_RD_PARITY   : in     vl_logic_vector(0 to 3);
        DMA_RD_DATA     : in     vl_logic_vector(0 to 31);
        CS1             : in     vl_logic;
        CS0_N           : in     vl_logic;
        CODE7           : in     vl_logic_vector(7 downto 0);
        CODE6           : in     vl_logic_vector(7 downto 0);
        CODE5           : in     vl_logic_vector(7 downto 0);
        CODE4           : in     vl_logic_vector(7 downto 0);
        CODE3           : in     vl_logic_vector(7 downto 0);
        CODE2           : in     vl_logic_vector(7 downto 0);
        CODE1           : in     vl_logic_vector(7 downto 0);
        CODE0           : in     vl_logic_vector(7 downto 0);
        CHIPID          : in     vl_logic_vector(7 downto 0);
        CFG_RESET_N     : in     vl_logic;
        CFG_PRGM_N      : in     vl_logic;
        CFG_OSC         : in     vl_logic;
        CCLKIN          : in     vl_logic;
        BSRSO           : in     vl_logic;
        ADDR_HIGH_DEL_N : in     vl_logic;
        LPCS_INT        : in     vl_logic_vector(3 downto 0);
        RPCS_INT        : in     vl_logic_vector(3 downto 0)
    );
end sys_bus_top;
