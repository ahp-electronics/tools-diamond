library verilog;
use verilog.vl_types.all;
entity pmu_ctrl is
    generic(
        PMU_NPART       : integer := 1;
        PMUFSMTMR       : integer := 1;
        PMUCREGTMR      : integer := 1;
        PMUST_IDLE      : vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        PMUST_NORM      : vl_logic_vector(0 to 2) := (Hi0, Hi1, Hi1);
        PMUST_LPWR      : vl_logic_vector(0 to 2) := (Hi0, Hi1, Hi0);
        PMUST_STBY      : vl_logic_vector(0 to 2) := (Hi1, Hi0, Hi0);
        PMUST_SSLP      : vl_logic_vector(0 to 2) := (Hi1, Hi0, Hi1);
        PMUST_DSLP      : vl_logic_vector(0 to 2) := (Hi1, Hi1, Hi1);
        SEQST_IDLE      : vl_logic_vector(0 to 1) := (Hi0, Hi0);
        SEQST_ACT1      : vl_logic_vector(0 to 1) := (Hi1, Hi0);
        SEQST_ACT2      : vl_logic_vector(0 to 1) := (Hi1, Hi1);
        SEQST_ACT3      : vl_logic_vector(0 to 1) := (Hi0, Hi1)
    );
    port(
        pmu_uclk_sel    : out    vl_logic;
        pmu_lclk_dis    : out    vl_logic;
        pmu_cfgclk_en   : out    vl_logic;
        pmu_cfgpwr_en   : out    vl_logic;
        pmuwdtcnt_sel   : out    vl_logic_vector(1 downto 0);
        pmuwdt_set      : out    vl_logic;
        pmuwdt_run      : out    vl_logic;
        uwdt_start_ack  : out    vl_logic;
        pmu_uwdt_inten  : out    vl_logic;
        pmu_wdt_done    : out    vl_logic;
        pmu_refresh     : out    vl_logic;
        pmu_pseq_run    : out    vl_logic;
        pmu_psave_state : out    vl_logic;
        pmu_idle        : out    vl_logic;
        pmu_norm        : out    vl_logic;
        pmu_lpwr        : out    vl_logic;
        pmu_stby        : out    vl_logic;
        pmu_sslp        : out    vl_logic;
        pmu_dslp        : out    vl_logic;
        pmu_int_extpen  : out    vl_logic;
        pmu_int_sspien  : out    vl_logic;
        pmu_int_si2cen  : out    vl_logic;
        pmu_ip_en       : out    vl_logic;
        pmu_uwdt_en     : out    vl_logic;
        pmu_rst_async   : in     vl_logic;
        pmu_clk         : in     vl_logic;
        clk_dis_sense   : in     vl_logic;
        pmucr           : in     vl_logic_vector(7 downto 0);
        pmuwdtcr0       : in     vl_logic_vector(7 downto 0);
        pmuwdtcr1       : in     vl_logic_vector(7 downto 0);
        pmuwdt_fin      : in     vl_logic;
        pmuwdt_fin_m1   : in     vl_logic;
        mcr_uclk_sel    : in     vl_logic;
        programn_sync   : in     vl_logic;
        cfg_umode_sync  : in     vl_logic;
        cfg_pseq_busy_sync: in     vl_logic;
        cfg_pmu_int_sel_sync: in     vl_logic_vector(1 downto 0);
        cfg_pmu_int_sync: in     vl_logic;
        spiint_sync     : in     vl_logic;
        i2cint_sync     : in     vl_logic;
        extint_sync     : in     vl_logic;
        cibint_sel_sync : in     vl_logic_vector(1 downto 0);
        cibint_sync     : in     vl_logic;
        uwdt_start_set_sync: in     vl_logic;
        pmu_uwdt_en_sync: in     vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of PMU_NPART : constant is 1;
    attribute mti_svvh_generic_type of PMUFSMTMR : constant is 1;
    attribute mti_svvh_generic_type of PMUCREGTMR : constant is 1;
    attribute mti_svvh_generic_type of PMUST_IDLE : constant is 1;
    attribute mti_svvh_generic_type of PMUST_NORM : constant is 1;
    attribute mti_svvh_generic_type of PMUST_LPWR : constant is 1;
    attribute mti_svvh_generic_type of PMUST_STBY : constant is 1;
    attribute mti_svvh_generic_type of PMUST_SSLP : constant is 1;
    attribute mti_svvh_generic_type of PMUST_DSLP : constant is 1;
    attribute mti_svvh_generic_type of SEQST_IDLE : constant is 1;
    attribute mti_svvh_generic_type of SEQST_ACT1 : constant is 1;
    attribute mti_svvh_generic_type of SEQST_ACT2 : constant is 1;
    attribute mti_svvh_generic_type of SEQST_ACT3 : constant is 1;
end pmu_ctrl;
