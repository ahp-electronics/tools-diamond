library verilog;
use verilog.vl_types.all;
entity cfg_reg is
    generic(
        MASTER_SERI     : integer := 8;
        MASTER_PARA     : integer := 12;
        ASYNC_PERI      : integer := 13;
        SLAVE_SERI      : integer := 15;
        SLAVE_PARA      : integer := 9;
        FPSC_PARA       : integer := 7;
        MASTER_BYTE     : integer := 6;
        FLASH_SPI03     : integer := 5;
        FLASH_SPIX      : integer := 4;
        MPC_BYTE        : integer := 10;
        MPC_HWORD       : integer := 11;
        MPC_WORD        : integer := 14;
        CHK_PRE         : integer := 0;
        CHK_ID          : integer := 1;
        CHK_HDR         : integer := 2;
        CHK_FPGA        : integer := 3;
        CHK_RAM         : integer := 6;
        CHK_FPSC        : integer := 5;
        CHK_POST        : integer := 7;
        BUF_SIZE        : integer := 96;
        ADDR_WAIT0      : integer := 0;
        ADDR_WAIT1      : integer := 3;
        ADDR_WAIT2      : integer := 7;
        ADDR_LOAD       : integer := 2;
        ADDR_INCR       : integer := 4;
        ADDR_SHIFT      : integer := 6
    );
    port(
        SED_RDBK        : in     vl_logic;
        CCLK            : in     vl_logic;
        CFRONT_INIT_N   : in     vl_logic;
        LMODE           : in     vl_logic_vector(3 downto 0);
        DONE            : in     vl_logic;
        FSM_INIT_RAM    : in     vl_logic;
        FSM_RES_N       : in     vl_logic;
        CLR_WR_EN       : in     vl_logic;
        LAST_ADDR       : in     vl_logic_vector(13 downto 0);
        PARTID          : in     vl_logic_vector(31 downto 12);
        RD_CFG          : in     vl_logic;
        PRGM_JTAG       : in     vl_logic;
        PRGM_JTAG_N     : in     vl_logic;
        RD_CFG_JTAG     : in     vl_logic;
        TDI_JTAG        : in     vl_logic;
        RDBK_REG_RAM    : in     vl_logic;
        EN_CAPTURE_RAM  : in     vl_logic;
        EN_ONCE_RAM     : in     vl_logic;
        EN_RDBK_RAM     : in     vl_logic;
        EN_READCAP_RAM  : in     vl_logic;
        CAPT_I_N        : in     vl_logic;
        SYS_RD_CFG      : in     vl_logic;
        SYS_BUS_CFG     : in     vl_logic;
        SYS_DAISY       : in     vl_logic;
        RDBK_ADDR       : in     vl_logic_vector(13 downto 0);
        REPEAT_RDBK     : in     vl_logic;
        SYS_MODE        : in     vl_logic;
        EN_ADDR         : in     vl_logic;
        RDBK_PC_EN      : in     vl_logic;
        RDBK_ZERO_ALL_N : in     vl_logic;
        RDBK_DOUT       : in     vl_logic_vector(7 downto 0);
        DEL_D_REG       : in     vl_logic_vector(7 downto 0);
        P2S_REG0        : in     vl_logic;
        MASTER_SERI_DEC_REG: in     vl_logic;
        SYS_BUS_DEC     : in     vl_logic;
        SYS_RDBK        : out    vl_logic;
        READ_START      : out    vl_logic;
        CHK_STATE       : out    vl_logic_vector(2 downto 0);
        RAM_BIT_ERR     : out    vl_logic;
        FPSC_BIT_ERR    : out    vl_logic;
        RDBK_ADDR_ERR   : out    vl_logic;
        RST_ADDR_REG    : out    vl_logic;
        GOT_ADDR        : out    vl_logic;
        EN_ADDR_INCR    : out    vl_logic;
        SHIFT_ADDR_1ST  : out    vl_logic;
        SHIFT_ADDR_2ND  : out    vl_logic;
        BAD_ADDR        : out    vl_logic;
        GOT_DHEADER     : out    vl_logic;
        ERR_FLAG        : out    vl_logic_vector(1 downto 0);
        RST_DATA_REG_N  : in     vl_logic;
        GOT_DATA        : out    vl_logic;
        INIT_1_DATA     : out    vl_logic;
        SERIAL_DATA     : out    vl_logic;
        LD_RDBKD        : out    vl_logic;
        CFG_DATA        : out    vl_logic_vector(7 downto 0);
        RDBK_DATA       : out    vl_logic;
        RDBK_TDO_EN     : out    vl_logic;
        CAPTURE         : out    vl_logic;
        SYS_RDBKD       : out    vl_logic_vector(7 downto 0);
        RD_SHIFT        : out    vl_logic_vector(1 downto 0);
        RAMD_RDY        : out    vl_logic;
        RAMA_RDY        : out    vl_logic;
        FPSCD_RDY       : out    vl_logic;
        FPSCA_RDY       : out    vl_logic;
        SYS_BUSD        : out    vl_logic_vector(71 downto 0);
        SYS_BUSA        : out    vl_logic_vector(9 downto 0);
        MATCH           : out    vl_logic;
        ZERO_ALL_N      : out    vl_logic;
        GOT_POST        : out    vl_logic;
        IDCODE3         : out    vl_logic_vector(7 downto 0);
        IDCODE4         : out    vl_logic_vector(7 downto 0);
        IDCODE5         : out    vl_logic_vector(7 downto 0);
        IDCODE6         : out    vl_logic_vector(7 downto 0);
        IDCODE7         : out    vl_logic_vector(7 downto 0);
        DEC_EN          : out    vl_logic;
        OSC_SEL         : out    vl_logic_vector(2 downto 0)
    );
end cfg_reg;
