-- $Header: //synplicity/map202003lat/mappers/cpld/lib/gen_mach/dec.vhd#1 $
@ER--7R B:FRl8CkDRMoCC0sNFVsRHRDCVRFs#CkbsFOFDN5D0O0HC#RHbBvq]j6jj2vX
H
DLssN$ RQ 
 ;kR#CQ   38#0_oDFH4O_43ncN;DD
C

M00H$ R7B#RH
C
oMHCsOR5M:MRH0CCosU:=2
;
b0Fs5q

RH:RM0R#8F_Do_HOP0COFMs5-84RF0IMF2Rj;1

RF:Rk#0R0D8_FOoH_OPC05FsMR-48MFI0jFR22

;C

M78R 
B;
ONsECH0Os0kCeRp_B7 RRFV7R BH
#
ObFlFMMC0BReBR
RRsbF0R5
RRRRRRXRRRRRRRRRRRRRRRRRRRRRRRRRRRRR:FRRkR0RR71a_tpmQ:BR=4R''
2;CRM8ObFlFMMC0
;
ObFlFMMC0hRt7R
RRsbF0R5
RRRRRRXRRRRRRRRRRRRRRRRRRRRRRRRRRRRR:FRRkR0RR71a_tpmQ:BR=jR''
2;CRM8ObFlFMMC0
;
ObFlFMMC0BRBzz_1AR
RRsbF0R5
RRRRRRqjRRRRRRRRRRRRRRRRRRRRRRRRRRRR:HRRMRRRR71a_tpmQ
B;RRRRRjRARRRRRRRRRRRRRRRRRRRRRRRRRRRRRR:RHRMRRaR17m_pt;QB
RRRRBRRQRhRRRRRRRRRRRRRRRRRRRRRRRRRRRR:RRHMR1RRap7_mBtQ;R
RRRRR1RjRRRRRRRRRRRRRRRRRRRRRRRRRR:RRRkRF0RRR1_a7pQmtBR;
RRRRRzBmaRRRRRRRRRRRRRRRRRRRRRRRRRRR:FRRkR0RR71a_tpmQ;B2
8CMRlOFbCFMM
0;
H
#oDMNRsONsR$RR#:R0D8_FOoH_OPC05FsR4M-RI8FMR0Fj;R2
o#HMRNDO#FM0R_4:0R#8F_Do;HO
o#HMRNDO#FM0R_j:0R#8F_Do;HO
C
Lo
HMRRRRRRRRzR4:eRBBuam)Ruvq5=RX>FROM_#04
2;RRRRRRRRzR.:tRh7uam)RuvqRR5X=O>RF0M#_;j2
RRRRRRRR:zdRzBB_A1zR)umaqRvuq5R5,j2RMOF#40_,FROM_#041,R5,j2RsONsj$52
2;RRRRRRRRzRc:VRFsHMRHR04RF-RM4CRoMNCs0RC
RRRRRRRRRRRRRzRR.4_pRB:RB1z_zuARmR)av5quRHq52O,RF0M#_Rj,OsNs$-5H4R2,125H,NROs5s$H;22
RRRRRRRR8CMRMoCC0sNC
;
CRM8p7e_ 
B;




