library verilog;
use verilog.vl_types.all;
entity qd_spare_gate is
    port(
        signal_in       : in     vl_logic
    );
end qd_spare_gate;
