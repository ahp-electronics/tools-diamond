library verilog;
use verilog.vl_types.all;
entity BUFX16 is
    port(
        z               : out    vl_logic;
        a               : in     vl_logic
    );
end BUFX16;
