library verilog;
use verilog.vl_types.all;
entity DELC0P1 is
    port(
        A               : in     vl_logic;
        Z               : out    vl_logic
    );
end DELC0P1;
