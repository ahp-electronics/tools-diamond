library verilog;
use verilog.vl_types.all;
entity flash_block is
    port(
        fail_flash_a    : out    vl_logic;
        row_a           : out    vl_logic_vector(14 downto 0);
        ufm_row_sel_all_a: out    vl_logic;
        ufm_row_sel_none_a: out    vl_logic;
        cfg_row_sel_all_a: out    vl_logic;
        cfg_row_sel_none_a: out    vl_logic;
        trim_row_sel_all_a: out    vl_logic;
        trim_row_sel_none_a: out    vl_logic;
        feat_row_sel_all_a: out    vl_logic;
        feat_row_sel_none_a: out    vl_logic;
        subrow_mvena_ufm_a: out    vl_logic;
        subrow_mvenall_ufm_a: out    vl_logic;
        subrow_hvena_ufm_a: out    vl_logic;
        subrow_hvenall_ufm_a: out    vl_logic;
        subrow_mvena_cfg_a: out    vl_logic;
        subrow_mvenall_cfg_a: out    vl_logic;
        subrow_hvena_cfg_a: out    vl_logic;
        subrow_hvenall_cfg_a: out    vl_logic;
        subrow_mvena_tf_a: out    vl_logic;
        subrow_hvena_tf_a: out    vl_logic;
        sa_enall_a      : out    vl_logic;
        sa_ena_a        : out    vl_logic;
        wor_eval_a      : out    vl_logic;
        wand_eval_a     : out    vl_logic;
        era_ufm_a       : out    vl_logic;
        era_cfg_a       : out    vl_logic;
        era_trim_a      : out    vl_logic;
        era_feat_a      : out    vl_logic;
        prg_ufm_a       : out    vl_logic;
        prg_cfg_a       : out    vl_logic;
        prg_tf_a        : out    vl_logic;
        read_ufm_a      : out    vl_logic;
        read_cfg_a      : out    vl_logic;
        read_tf_a       : out    vl_logic;
        era_ver_a       : out    vl_logic;
        scp_a           : out    vl_logic;
        scpv_a          : out    vl_logic;
        softprg_a       : out    vl_logic;
        verify_a        : out    vl_logic;
        flash_en_a      : out    vl_logic;
        reg_enable_a    : out    vl_logic;
        sel_6p5v_a      : out    vl_logic;
        fl_ready_rst_a  : out    vl_logic;
        fl_erase_cfg0   : out    vl_logic;
        fl_erase_ufm0   : out    vl_logic;
        fl_erase_trim   : out    vl_logic;
        fl_erase_fea    : out    vl_logic;
        mux32_out1_a    : out    vl_logic;
        mux32_out2_a    : out    vl_logic;
        pwtc_well_a     : out    vl_logic;
        erase_setup_a   : out    vl_logic;
        erase_pulse_a   : out    vl_logic;
        erapdis_a       : out    vl_logic;
        prg_pwtc_a      : out    vl_logic;
        prog_disch_a    : out    vl_logic;
        en_vreg_mon_a   : out    vl_logic;
        prgdrv_ena_a    : out    vl_logic;
        col_shift_a     : out    vl_logic;
        colstart_a      : out    vl_logic_vector(3 downto 0);
        col_rst_a       : out    vl_logic;
        readpart_a      : out    vl_logic_vector(3 downto 0);
        capture_dout_a  : out    vl_logic;
        src_clamp_a     : out    vl_logic;
        drain_ctrl_a    : out    vl_logic;
        prestep_in_neg_a: out    vl_logic_vector(2 downto 0);
        step_in_neg_a   : out    vl_logic_vector(2 downto 0);
        prg_pulse_a     : out    vl_logic_vector(3 downto 0);
        prgdrv_enall_a  : out    vl_logic;
        ppt_en_a        : out    vl_logic;
        ppt_rowsel_a    : out    vl_logic;
        ppt_pset_a      : out    vl_logic;
        fl_load_trim0   : out    vl_logic;
        fl_load_trim1   : out    vl_logic;
        fl_load_pes     : out    vl_logic;
        fl_load_mes     : out    vl_logic;
        fl_load_uds_trn : out    vl_logic;
        fl_load_tss     : out    vl_logic;
        fl_load_pwd     : out    vl_logic;
        fl_load_fea     : out    vl_logic;
        fl_load_feabits : out    vl_logic;
        fl_load_fss     : out    vl_logic;
        fl_load_udss0   : out    vl_logic;
        fl_load_ufs0    : out    vl_logic;
        device_a        : in     vl_logic_vector(2 downto 0);
        l_row_cfg_a     : in     vl_logic;
        l_row_ufm_a     : in     vl_logic;
        fl_dout_a       : in     vl_logic_vector(63 downto 0);
        fl_ready_a      : in     vl_logic;
        vwlp_active_a   : in     vl_logic;
        neg_edge_det_a  : in     vl_logic;
        well_active_a   : in     vl_logic;
        ready_vfy_a     : in     vl_logic;
        c_bl_a          : in     vl_logic_vector(3 downto 0);
        lastcol_a       : in     vl_logic_vector(3 downto 0);
        fail_flash_b    : out    vl_logic;
        row_b           : out    vl_logic_vector(14 downto 0);
        ufm_row_sel_all_b: out    vl_logic;
        ufm_row_sel_none_b: out    vl_logic;
        cfg_row_sel_all_b: out    vl_logic;
        cfg_row_sel_none_b: out    vl_logic;
        trim_row_sel_all_b: out    vl_logic;
        trim_row_sel_none_b: out    vl_logic;
        feat_row_sel_all_b: out    vl_logic;
        feat_row_sel_none_b: out    vl_logic;
        subrow_mvena_ufm_b: out    vl_logic;
        subrow_mvenall_ufm_b: out    vl_logic;
        subrow_hvena_ufm_b: out    vl_logic;
        subrow_hvenall_ufm_b: out    vl_logic;
        subrow_mvena_cfg_b: out    vl_logic;
        subrow_mvenall_cfg_b: out    vl_logic;
        subrow_hvena_cfg_b: out    vl_logic;
        subrow_hvenall_cfg_b: out    vl_logic;
        subrow_mvena_tf_b: out    vl_logic;
        subrow_hvena_tf_b: out    vl_logic;
        sa_enall_b      : out    vl_logic;
        sa_ena_b        : out    vl_logic;
        wor_eval_b      : out    vl_logic;
        wand_eval_b     : out    vl_logic;
        era_ufm_b       : out    vl_logic;
        era_cfg_b       : out    vl_logic;
        era_trim_b      : out    vl_logic;
        era_feat_b      : out    vl_logic;
        prg_ufm_b       : out    vl_logic;
        prg_cfg_b       : out    vl_logic;
        prg_tf_b        : out    vl_logic;
        read_ufm_b      : out    vl_logic;
        read_cfg_b      : out    vl_logic;
        read_tf_b       : out    vl_logic;
        era_ver_b       : out    vl_logic;
        scp_b           : out    vl_logic;
        scpv_b          : out    vl_logic;
        softprg_b       : out    vl_logic;
        verify_b        : out    vl_logic;
        flash_en_b      : out    vl_logic;
        reg_enable_b    : out    vl_logic;
        sel_6p5v_b      : out    vl_logic;
        fl_ready_rst_b  : out    vl_logic;
        fl_erase_cfg1   : out    vl_logic;
        fl_erase_ufm1   : out    vl_logic;
        fl_erase_pubkey : out    vl_logic;
        fl_erase_csec   : out    vl_logic;
        mux32_out1_b    : out    vl_logic;
        mux32_out2_b    : out    vl_logic;
        pwtc_well_b     : out    vl_logic;
        erase_setup_b   : out    vl_logic;
        erase_pulse_b   : out    vl_logic;
        erapdis_b       : out    vl_logic;
        prg_pwtc_b      : out    vl_logic;
        prog_disch_b    : out    vl_logic;
        en_vreg_mon_b   : out    vl_logic;
        prgdrv_ena_b    : out    vl_logic;
        col_shift_b     : out    vl_logic;
        colstart_b      : out    vl_logic_vector(3 downto 0);
        col_rst_b       : out    vl_logic;
        readpart_b      : out    vl_logic_vector(3 downto 0);
        capture_dout_b  : out    vl_logic;
        src_clamp_b     : out    vl_logic;
        drain_ctrl_b    : out    vl_logic;
        prestep_in_neg_b: out    vl_logic_vector(2 downto 0);
        step_in_neg_b   : out    vl_logic_vector(2 downto 0);
        prg_pulse_b     : out    vl_logic_vector(3 downto 0);
        prgdrv_enall_b  : out    vl_logic;
        ppt_en_b        : out    vl_logic;
        ppt_rowsel_b    : out    vl_logic;
        ppt_pset_b      : out    vl_logic;
        fl_load_pkey0   : out    vl_logic;
        fl_load_pkey1   : out    vl_logic;
        fl_load_pkey2   : out    vl_logic;
        fl_load_pkey3   : out    vl_logic;
        fl_load_csec    : out    vl_logic;
        fl_load_udss1   : out    vl_logic;
        fl_load_ufs1    : out    vl_logic;
        fl_load_pks     : out    vl_logic;
        fl_load_css     : out    vl_logic;
        device_b        : in     vl_logic_vector(2 downto 0);
        l_row_cfg_b     : in     vl_logic;
        l_row_ufm_b     : in     vl_logic;
        fl_dout_b       : in     vl_logic_vector(63 downto 0);
        fl_ready_b      : in     vl_logic;
        vwlp_active_b   : in     vl_logic;
        neg_edge_det_b  : in     vl_logic;
        well_active_b   : in     vl_logic;
        ready_vfy_b     : in     vl_logic;
        c_bl_b          : in     vl_logic_vector(3 downto 0);
        lastcol_b       : in     vl_logic_vector(3 downto 0);
        fail_flash_c    : out    vl_logic;
        row_c           : out    vl_logic_vector(14 downto 0);
        ufm_row_sel_all_c: out    vl_logic;
        ufm_row_sel_none_c: out    vl_logic;
        cfg_row_sel_all_c: out    vl_logic;
        cfg_row_sel_none_c: out    vl_logic;
        trim_row_sel_all_c: out    vl_logic;
        trim_row_sel_none_c: out    vl_logic;
        feat_row_sel_all_c: out    vl_logic;
        feat_row_sel_none_c: out    vl_logic;
        subrow_mvena_ufm_c: out    vl_logic;
        subrow_mvenall_ufm_c: out    vl_logic;
        subrow_hvena_ufm_c: out    vl_logic;
        subrow_hvenall_ufm_c: out    vl_logic;
        subrow_mvena_cfg_c: out    vl_logic;
        subrow_mvenall_cfg_c: out    vl_logic;
        subrow_hvena_cfg_c: out    vl_logic;
        subrow_hvenall_cfg_c: out    vl_logic;
        subrow_mvena_tf_c: out    vl_logic;
        subrow_hvena_tf_c: out    vl_logic;
        sa_enall_c      : out    vl_logic;
        sa_ena_c        : out    vl_logic;
        wor_eval_c      : out    vl_logic;
        wand_eval_c     : out    vl_logic;
        era_ufm_c       : out    vl_logic;
        era_cfg_c       : out    vl_logic;
        era_trim_c      : out    vl_logic;
        era_feat_c      : out    vl_logic;
        prg_ufm_c       : out    vl_logic;
        prg_cfg_c       : out    vl_logic;
        prg_tf_c        : out    vl_logic;
        read_ufm_c      : out    vl_logic;
        read_cfg_c      : out    vl_logic;
        read_tf_c       : out    vl_logic;
        era_ver_c       : out    vl_logic;
        scp_c           : out    vl_logic;
        scpv_c          : out    vl_logic;
        softprg_c       : out    vl_logic;
        verify_c        : out    vl_logic;
        flash_en_c      : out    vl_logic;
        reg_enable_c    : out    vl_logic;
        sel_6p5v_c      : out    vl_logic;
        fl_ready_rst_c  : out    vl_logic;
        fl_erase_ufm2   : out    vl_logic;
        fl_erase_ufm3   : out    vl_logic;
        fl_erase_aeskey : out    vl_logic;
        fl_erase_usec   : out    vl_logic;
        mux32_out1_c    : out    vl_logic;
        mux32_out2_c    : out    vl_logic;
        pwtc_well_c     : out    vl_logic;
        erase_setup_c   : out    vl_logic;
        erase_pulse_c   : out    vl_logic;
        erapdis_c       : out    vl_logic;
        prg_pwtc_c      : out    vl_logic;
        prog_disch_c    : out    vl_logic;
        en_vreg_mon_c   : out    vl_logic;
        prgdrv_ena_c    : out    vl_logic;
        col_shift_c     : out    vl_logic;
        colstart_c      : out    vl_logic_vector(3 downto 0);
        col_rst_c       : out    vl_logic;
        readpart_c      : out    vl_logic_vector(3 downto 0);
        capture_dout_c  : out    vl_logic;
        src_clamp_c     : out    vl_logic;
        drain_ctrl_c    : out    vl_logic;
        prestep_in_neg_c: out    vl_logic_vector(2 downto 0);
        step_in_neg_c   : out    vl_logic_vector(2 downto 0);
        prg_pulse_c     : out    vl_logic_vector(3 downto 0);
        prgdrv_enall_c  : out    vl_logic;
        ppt_en_c        : out    vl_logic;
        ppt_rowsel_c    : out    vl_logic;
        ppt_pset_c      : out    vl_logic;
        fl_load_akey0   : out    vl_logic;
        fl_load_akey1   : out    vl_logic;
        fl_load_usec    : out    vl_logic;
        fl_load_ufs2    : out    vl_logic;
        fl_load_ufs3    : out    vl_logic;
        fl_load_aks     : out    vl_logic;
        fl_load_uss     : out    vl_logic;
        device_c        : in     vl_logic_vector(2 downto 0);
        l_row_cfg_c     : in     vl_logic;
        l_row_ufm_c     : in     vl_logic;
        fl_dout_c       : in     vl_logic_vector(63 downto 0);
        fl_ready_c      : in     vl_logic;
        vwlp_active_c   : in     vl_logic;
        neg_edge_det_c  : in     vl_logic;
        well_active_c   : in     vl_logic;
        ready_vfy_c     : in     vl_logic;
        c_bl_c          : in     vl_logic_vector(3 downto 0);
        lastcol_c       : in     vl_logic_vector(3 downto 0);
        fail_flash      : out    vl_logic;
        flash_clk_mfg   : out    vl_logic;
        fl_modal_state  : out    vl_logic_vector(31 downto 0);
        fl_er_count     : out    vl_logic_vector(11 downto 0);
        fl_pg_count     : out    vl_logic_vector(9 downto 0);
        lsc_sdm         : out    vl_logic;
        lsc_sdm_cfg0    : out    vl_logic;
        lsc_sdm_cfg1    : out    vl_logic;
        fl_finish_ppt   : out    vl_logic;
        fl_busy_ppt     : out    vl_logic;
        ppt_init_tsf_asr_exec: out    vl_logic;
        ppt_write_incr_exec: out    vl_logic;
        ppt_dat         : out    vl_logic_vector(7 downto 0);
        ppt_dsr_shf8_en : out    vl_logic;
        ppt_dsr_shf     : out    vl_logic;
        fl_finish_cdm   : out    vl_logic;
        fl_busy_cdm     : out    vl_logic;
        fl_finish_sdm   : out    vl_logic;
        fl_busy_sdm     : out    vl_logic;
        fail_sdm_a      : out    vl_logic;
        fail_sdm_b      : out    vl_logic;
        sdm_start_bse   : out    vl_logic;
        sdm_bse_eof     : out    vl_logic;
        preamble_std_sdm: out    vl_logic;
        preamble_enc_sdm: out    vl_logic;
        preamble_err_sdm: out    vl_logic;
        sdm_init_sram_asr_exec: out    vl_logic;
        dnld_dat        : out    vl_logic_vector(7 downto 0);
        dnld_dat_en     : out    vl_logic;
        ppt_fail        : out    vl_logic;
        por             : in     vl_logic;
        isc_rst_async   : in     vl_logic;
        isc_rst_sync    : in     vl_logic;
        smclk           : in     vl_logic;
        fl_smclk_mfg    : in     vl_logic;
        scanen          : in     vl_logic;
        isc_exec_a      : in     vl_logic;
        isc_exec_b      : in     vl_logic;
        isc_exec_c      : in     vl_logic;
        isc_exec_d      : in     vl_logic;
        isc_exec_e      : in     vl_logic;
        mfg_margin_en   : in     vl_logic;
        mfg_skip_era    : in     vl_logic;
        mfg_skip_ev     : in     vl_logic;
        mfg_skip_prgvfy : in     vl_logic;
        mfg_skip_scp    : in     vl_logic;
        mfg_skip_softprg: in     vl_logic;
        mfg_vreg_mon    : in     vl_logic;
        mfg_nofail      : in     vl_logic;
        mfg_dis_sel6p5v : in     vl_logic;
        mfg_4xprg       : in     vl_logic;
        mfg_step_size   : in     vl_logic;
        mfg_ers_cnt     : in     vl_logic_vector(3 downto 0);
        mfg_ers_perstep : in     vl_logic_vector(1 downto 0);
        mfg_ers_steps   : in     vl_logic_vector(1 downto 0);
        mfg_prg_cnt     : in     vl_logic_vector(2 downto 0);
        mfg_sp_cnt      : in     vl_logic_vector(2 downto 0);
        mfg_scp_cnt     : in     vl_logic_vector(2 downto 0);
        mfg_fl_enable   : in     vl_logic;
        mfg_mux1_sel    : in     vl_logic_vector(4 downto 0);
        mfg_mux2_sel    : in     vl_logic_vector(4 downto 0);
        mfg_fl_sel      : in     vl_logic_vector(1 downto 0);
        mfg_fl_pe       : in     vl_logic;
        mfg_fl_pp       : in     vl_logic;
        mfg_mtest_fl_sel: in     vl_logic_vector(1 downto 0);
        trim_row_ev     : in     vl_logic;
        trim_sel6p5v    : in     vl_logic;
        trim_ers_pw     : in     vl_logic_vector(2 downto 0);
        trim_prg_pw     : in     vl_logic_vector(2 downto 0);
        trim_scp_pw     : in     vl_logic_vector(2 downto 0);
        trim_verify     : in     vl_logic_vector(1 downto 0);
        trim_neg_init_a : in     vl_logic_vector(5 downto 0);
        trim_neg_init_b : in     vl_logic_vector(5 downto 0);
        trim_neg_init_c : in     vl_logic_vector(5 downto 0);
        trim_fl_pe_en   : in     vl_logic;
        access_flash_all: in     vl_logic;
        fsafe           : in     vl_logic;
        mfg_ppt_abort   : in     vl_logic;
        fl_start_ppt    : in     vl_logic;
        fl_start_cdm    : in     vl_logic;
        fl_start_sdm_cfg0: in     vl_logic;
        fl_start_sdm_cfg1: in     vl_logic;
        authdone_sdm0_start: in     vl_logic;
        authdone_sdm1_start: in     vl_logic;
        dev_sdm_cfg0_exec: in     vl_logic;
        dev_sdm_cfg1_exec: in     vl_logic;
        busy_sram       : in     vl_logic;
        finish_bse      : in     vl_logic;
        fail_bse        : in     vl_logic;
        njbse_preamble  : in     vl_logic;
        sdm_run         : in     vl_logic;
        mc1_ppt_bits    : in     vl_logic_vector(7 downto 0);
        busy_flash      : out    vl_logic;
        fl_exec_buf     : out    vl_logic_vector(127 downto 0);
        current_sector  : out    vl_logic_vector(11 downto 0);
        mfg_flash_en    : in     vl_logic;
        access_sudo     : in     vl_logic;
        fl_erase_all_qual: in     vl_logic;
        fl_erase_qual   : in     vl_logic;
        fl_erase_exec   : in     vl_logic;
        fl_prog_ucode_qual: in     vl_logic;
        fl_prog_done_qual: in     vl_logic;
        fl_prog_sec_qual: in     vl_logic;
        fl_prog_secplus_qual: in     vl_logic;
        fl_disable_done0_qual: in     vl_logic;
        fl_disable_done1_qual: in     vl_logic;
        fl_udss0_authdone_exec: in     vl_logic;
        fl_udss1_authdone_exec: in     vl_logic;
        fl_prog_uds_qual: in     vl_logic;
        fl_prog_authmode_qual: in     vl_logic;
        fl_prog_aesfea_qual: in     vl_logic;
        fl_init_addr_qual: in     vl_logic;
        fl_write_addr_qual: in     vl_logic;
        fl_prog_incr_nv_qual: in     vl_logic;
        fl_read_incr_nv_qual: in     vl_logic;
        fl_prog_password_qual: in     vl_logic;
        fl_prog_feature_qual: in     vl_logic;
        fl_prog_feabits_qual: in     vl_logic;
        fl_init_addr_ufm_qual: in     vl_logic;
        fl_prog_tag_qual: in     vl_logic;
        fl_erase_tag_qual: in     vl_logic;
        fl_read_tag_qual: in     vl_logic;
        fl_prog_pes_qual: in     vl_logic;
        fl_prog_mes_qual: in     vl_logic;
        fl_prog_hes_qual: in     vl_logic;
        fl_prog_trim0_qual: in     vl_logic;
        fl_prog_trim1_qual: in     vl_logic;
        fl_read_hes_qual: in     vl_logic;
        fl_mtest_qual   : in     vl_logic;
        fl_prog_pubkey0_qual: in     vl_logic;
        fl_prog_pubkey1_qual: in     vl_logic;
        fl_prog_pubkey2_qual: in     vl_logic;
        fl_prog_pubkey3_qual: in     vl_logic;
        fl_prog_aeskey0_qual: in     vl_logic;
        fl_prog_aeskey1_qual: in     vl_logic;
        fl_prog_usec_qual: in     vl_logic;
        fl_prog_csec_qual: in     vl_logic;
        buf128_dat      : in     vl_logic_vector(127 downto 0);
        sector_dat      : in     vl_logic_vector(15 downto 0);
        sector_erase    : in     vl_logic_vector(11 downto 0);
        ppt_timer_en    : in     vl_logic
    );
end flash_block;
