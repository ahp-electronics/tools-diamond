library verilog;
use verilog.vl_types.all;
entity i2c_port is
    generic(
        TR_IDLE         : vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        TR_ADDR         : vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi1);
        TR_ACKA         : vl_logic_vector(0 to 2) := (Hi0, Hi1, Hi1);
        TR_INFO         : vl_logic_vector(0 to 2) := (Hi0, Hi1, Hi0);
        TR_ACKB         : vl_logic_vector(0 to 2) := (Hi1, Hi1, Hi0);
        TR_RDAT         : vl_logic_vector(0 to 2) := (Hi1, Hi1, Hi1);
        TR_ACKD         : vl_logic_vector(0 to 2) := (Hi1, Hi0, Hi1);
        MC_IDLE         : vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi0);
        MC_STAP         : vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi1, Hi0);
        MC_STAA         : vl_logic_vector(0 to 3) := (Hi1, Hi0, Hi0, Hi0);
        MC_STAB         : vl_logic_vector(0 to 3) := (Hi1, Hi0, Hi0, Hi1);
        MC_STAC         : vl_logic_vector(0 to 3) := (Hi1, Hi0, Hi1, Hi1);
        MC_STAD         : vl_logic_vector(0 to 3) := (Hi1, Hi0, Hi1, Hi0);
        MC_TRCA         : vl_logic_vector(0 to 3) := (Hi1, Hi1, Hi1, Hi0);
        MC_TRCB         : vl_logic_vector(0 to 3) := (Hi1, Hi1, Hi1, Hi1);
        MC_TRCC         : vl_logic_vector(0 to 3) := (Hi1, Hi1, Hi0, Hi1);
        MC_TRCD         : vl_logic_vector(0 to 3) := (Hi1, Hi1, Hi0, Hi0);
        MC_STRP         : vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi1, Hi1);
        MC_STOP         : vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi1);
        MC_STOA         : vl_logic_vector(0 to 3) := (Hi0, Hi1, Hi0, Hi0);
        MC_STOB         : vl_logic_vector(0 to 3) := (Hi0, Hi1, Hi1, Hi0);
        MC_STOC         : vl_logic_vector(0 to 3) := (Hi0, Hi1, Hi1, Hi1);
        MC_STOD         : vl_logic_vector(0 to 3) := (Hi0, Hi1, Hi0, Hi1)
    );
    port(
        sda_out         : out    vl_logic;
        sda_oe          : out    vl_logic;
        scl_out         : out    vl_logic;
        scl_oe          : out    vl_logic;
        i2crxdr         : out    vl_logic_vector(7 downto 0);
        i2cgcdr         : out    vl_logic_vector(7 downto 0);
        i2csr           : out    vl_logic_vector(7 downto 0);
        i2c_hsmode      : out    vl_logic;
        i2c_wkup        : out    vl_logic;
        ADDR_LSB_USR    : in     vl_logic_vector(1 downto 0);
        i2c_rst_async   : in     vl_logic;
        sda_in          : in     vl_logic;
        scl_in          : in     vl_logic;
        del_clk         : in     vl_logic;
        sb_clk_i        : in     vl_logic;
        i2ccr1          : in     vl_logic_vector(7 downto 0);
        i2ccmdr         : in     vl_logic_vector(7 downto 0);
        i2ctxdr         : in     vl_logic_vector(7 downto 0);
        i2cbr           : in     vl_logic_vector(9 downto 0);
        i2csaddr        : in     vl_logic_vector(7 downto 0);
        i2ccr1_wt       : in     vl_logic;
        i2ccmdr_wt      : in     vl_logic;
        i2cbr_wt        : in     vl_logic;
        i2ctxdr_wt      : in     vl_logic;
        i2csaddr_wt     : in     vl_logic;
        i2crxdr_rd      : in     vl_logic;
        i2cgcdr_rd      : in     vl_logic;
        trim_sda_del    : in     vl_logic_vector(3 downto 0);
        scan_test_mode  : in     vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of TR_IDLE : constant is 1;
    attribute mti_svvh_generic_type of TR_ADDR : constant is 1;
    attribute mti_svvh_generic_type of TR_ACKA : constant is 1;
    attribute mti_svvh_generic_type of TR_INFO : constant is 1;
    attribute mti_svvh_generic_type of TR_ACKB : constant is 1;
    attribute mti_svvh_generic_type of TR_RDAT : constant is 1;
    attribute mti_svvh_generic_type of TR_ACKD : constant is 1;
    attribute mti_svvh_generic_type of MC_IDLE : constant is 1;
    attribute mti_svvh_generic_type of MC_STAP : constant is 1;
    attribute mti_svvh_generic_type of MC_STAA : constant is 1;
    attribute mti_svvh_generic_type of MC_STAB : constant is 1;
    attribute mti_svvh_generic_type of MC_STAC : constant is 1;
    attribute mti_svvh_generic_type of MC_STAD : constant is 1;
    attribute mti_svvh_generic_type of MC_TRCA : constant is 1;
    attribute mti_svvh_generic_type of MC_TRCB : constant is 1;
    attribute mti_svvh_generic_type of MC_TRCC : constant is 1;
    attribute mti_svvh_generic_type of MC_TRCD : constant is 1;
    attribute mti_svvh_generic_type of MC_STRP : constant is 1;
    attribute mti_svvh_generic_type of MC_STOP : constant is 1;
    attribute mti_svvh_generic_type of MC_STOA : constant is 1;
    attribute mti_svvh_generic_type of MC_STOB : constant is 1;
    attribute mti_svvh_generic_type of MC_STOC : constant is 1;
    attribute mti_svvh_generic_type of MC_STOD : constant is 1;
end i2c_port;
