library verilog;
use verilog.vl_types.all;
entity cfg_pdec is
    port(
        por             : in     vl_logic;
        smclk           : in     vl_logic;
        isc_done        : in     vl_logic;
        wkup_done       : in     vl_logic;
        ctrl_sspi_auto  : in     vl_logic;
        ctrl_cpu_manu   : in     vl_logic;
        cfg_pin         : in     vl_logic_vector(2 downto 0);
        programn_pin    : in     vl_logic;
        initn_pin       : in     vl_logic;
        done_pin        : in     vl_logic;
        gsrn_pin        : in     vl_logic;
        mspisel_pin     : in     vl_logic_vector(3 downto 0);
        sspi_csn        : in     vl_logic;
        scpu_csn        : in     vl_logic;
        csn_pin         : in     vl_logic_vector(1 downto 0);
        i2c_cfg_active  : in     vl_logic;
        wbc_cfg_active  : in     vl_logic;
        njboot_dat      : in     vl_logic_vector(7 downto 0);
        jtag_active_smsync_jb: in     vl_logic;
        mc1_persist_mspi: in     vl_logic;
        mc1_persist_sspi: in     vl_logic;
        mc1_persist_i2c : in     vl_logic;
        mc1_persist_cpu8: in     vl_logic;
        mc1_persist_cpu16: in     vl_logic;
        fsd_persistn_progn: in     vl_logic;
        fsd_persist_initn: in     vl_logic;
        fsd_persist_done: in     vl_logic;
        fsd_persist_mspi: in     vl_logic;
        fsd_persistn_sspi: in     vl_logic;
        fsd_persistn_i2c: in     vl_logic;
        fsd_boot_sel    : in     vl_logic_vector(2 downto 0);
        fifo_rst        : in     vl_logic;
        mfg_scpu_en     : in     vl_logic;
        cfg0_latter     : in     vl_logic;
        persist_mspi    : out    vl_logic;
        persist_sspi    : out    vl_logic;
        persist_i2c     : out    vl_logic;
        persist_cpu8    : out    vl_logic;
        persist_cpu16   : out    vl_logic;
        p_slave         : out    vl_logic;
        p_slave_manu    : out    vl_logic;
        p_mspi0         : out    vl_logic;
        p_mspim         : out    vl_logic;
        p_scm           : out    vl_logic;
        p_sspi          : out    vl_logic;
        p_sp8           : out    vl_logic;
        p_sp16          : out    vl_logic;
        p_i2c           : out    vl_logic;
        p_scpu          : out    vl_logic;
        p_mspi_slow     : out    vl_logic;
        p_mspi_fast     : out    vl_logic;
        p_mspi_dual     : out    vl_logic;
        p_mspi_quad     : out    vl_logic;
        p_mp8           : out    vl_logic;
        p_mp16          : out    vl_logic;
        p_mp8_quad      : out    vl_logic;
        p_mp16_quad     : out    vl_logic;
        p_sst           : out    vl_logic;
        p_mspi_all      : out    vl_logic;
        p_end_bpft      : out    vl_logic;
        njport_init     : out    vl_logic;
        njport_active   : out    vl_logic;
        njport_exec     : out    vl_logic;
        wbc_active      : out    vl_logic;
        sspi_active     : out    vl_logic;
        i2c_active      : out    vl_logic;
        p_eboot0p       : out    vl_logic;
        p_eboot1p       : out    vl_logic;
        p_eboot1s       : out    vl_logic;
        p_eboot2p       : out    vl_logic;
        p_eboot2s       : out    vl_logic;
        p_nboot         : out    vl_logic;
        p_iboot0p       : out    vl_logic;
        p_iboot1p       : out    vl_logic;
        p_iboot1s       : out    vl_logic;
        p_iboot2p       : out    vl_logic;
        p_iboot2s       : out    vl_logic;
        programn_tog    : out    vl_logic;
        programn_pin_sync: out    vl_logic;
        initn_pin_sync  : out    vl_logic;
        done_pin_sync   : out    vl_logic;
        done_rise1      : out    vl_logic;
        gsrn_pin_sync   : out    vl_logic;
        boot_setup      : out    vl_logic_vector(5 downto 0);
        persist_slave   : out    vl_logic;
        p_iboot0s       : out    vl_logic
    );
end cfg_pdec;
