library verilog;
use verilog.vl_types.all;
entity PCSA_sim is
    generic(
        CONFIG_FILE     : string  := "configfile.txt";
        BASE_ADDRESS    : string  := "0x36000"
    );
    port(
        HDINP0          : in     vl_logic;
        HDINN0          : in     vl_logic;
        HDINP1          : in     vl_logic;
        HDINN1          : in     vl_logic;
        HDINP2          : in     vl_logic;
        HDINN2          : in     vl_logic;
        HDINP3          : in     vl_logic;
        HDINN3          : in     vl_logic;
        REFCLKP         : in     vl_logic;
        REFCLKN         : in     vl_logic;
        RXREFCLKP       : in     vl_logic;
        RXREFCLKN       : in     vl_logic;
        HDOUTP0         : out    vl_logic;
        HDOUTN0         : out    vl_logic;
        HDOUTP1         : out    vl_logic;
        HDOUTN1         : out    vl_logic;
        HDOUTP2         : out    vl_logic;
        HDOUTN2         : out    vl_logic;
        HDOUTP3         : out    vl_logic;
        HDOUTN3         : out    vl_logic;
        FFC_QUAD_RST    : in     vl_logic;
        FFC_MACRO_RST   : in     vl_logic;
        FFC_LANE_TX_RST0: in     vl_logic;
        FFC_LANE_TX_RST1: in     vl_logic;
        FFC_LANE_TX_RST2: in     vl_logic;
        FFC_LANE_TX_RST3: in     vl_logic;
        FFC_LANE_RX_RST0: in     vl_logic;
        FFC_LANE_RX_RST1: in     vl_logic;
        FFC_LANE_RX_RST2: in     vl_logic;
        FFC_LANE_RX_RST3: in     vl_logic;
        FFC_PCIE_EI_EN_0: in     vl_logic;
        FFC_PCIE_EI_EN_1: in     vl_logic;
        FFC_PCIE_EI_EN_2: in     vl_logic;
        FFC_PCIE_EI_EN_3: in     vl_logic;
        FFC_PCIE_CT_0   : in     vl_logic;
        FFC_PCIE_CT_1   : in     vl_logic;
        FFC_PCIE_CT_2   : in     vl_logic;
        FFC_PCIE_CT_3   : in     vl_logic;
        FFC_PCIE_TX_0   : in     vl_logic;
        FFC_PCIE_TX_1   : in     vl_logic;
        FFC_PCIE_TX_2   : in     vl_logic;
        FFC_PCIE_TX_3   : in     vl_logic;
        FFC_PCIE_RX_0   : in     vl_logic;
        FFC_PCIE_RX_1   : in     vl_logic;
        FFC_PCIE_RX_2   : in     vl_logic;
        FFC_PCIE_RX_3   : in     vl_logic;
        FFC_SD_0        : in     vl_logic;
        FFC_SD_1        : in     vl_logic;
        FFC_SD_2        : in     vl_logic;
        FFC_SD_3        : in     vl_logic;
        FFC_EN_CGA_0    : in     vl_logic;
        FFC_EN_CGA_1    : in     vl_logic;
        FFC_EN_CGA_2    : in     vl_logic;
        FFC_EN_CGA_3    : in     vl_logic;
        FFC_ALIGN_EN_0  : in     vl_logic;
        FFC_ALIGN_EN_1  : in     vl_logic;
        FFC_ALIGN_EN_2  : in     vl_logic;
        FFC_ALIGN_EN_3  : in     vl_logic;
        FFC_AB_RESET    : in     vl_logic;
        FFC_CD_RESET    : in     vl_logic;
        FFC_FB_LB_0     : in     vl_logic;
        FFC_FB_LB_1     : in     vl_logic;
        FFC_FB_LB_2     : in     vl_logic;
        FFC_FB_LB_3     : in     vl_logic;
        FFC_SB_INV_RX_0 : in     vl_logic;
        FFC_SB_INV_RX_1 : in     vl_logic;
        FFC_SB_INV_RX_2 : in     vl_logic;
        FFC_SB_INV_RX_3 : in     vl_logic;
        FFS_PCIE_CON_0  : out    vl_logic;
        FFS_PCIE_CON_1  : out    vl_logic;
        FFS_PCIE_CON_2  : out    vl_logic;
        FFS_PCIE_CON_3  : out    vl_logic;
        FFS_PCIE_DONE_0 : out    vl_logic;
        FFS_PCIE_DONE_1 : out    vl_logic;
        FFS_PCIE_DONE_2 : out    vl_logic;
        FFS_PCIE_DONE_3 : out    vl_logic;
        FFS_LS_STATUS_0 : out    vl_logic;
        FFS_LS_STATUS_1 : out    vl_logic;
        FFS_LS_STATUS_2 : out    vl_logic;
        FFS_LS_STATUS_3 : out    vl_logic;
        FFS_AB_STATUS   : out    vl_logic;
        FFS_CD_STATUS   : out    vl_logic;
        FFS_AB_ALIGNED  : out    vl_logic;
        FFS_CD_ALIGNED  : out    vl_logic;
        FFS_AB_FAILED   : out    vl_logic;
        FFS_CD_FAILED   : out    vl_logic;
        FFS_CC_ORUN_0   : out    vl_logic;
        FFS_CC_ORUN_1   : out    vl_logic;
        FFS_CC_ORUN_2   : out    vl_logic;
        FFS_CC_ORUN_3   : out    vl_logic;
        FFS_CC_URUN_0   : out    vl_logic;
        FFS_CC_URUN_1   : out    vl_logic;
        FFS_CC_URUN_2   : out    vl_logic;
        FFS_CC_URUN_3   : out    vl_logic;
        FFS_RLOS_LO0    : out    vl_logic;
        FFS_RLOS_LO1    : out    vl_logic;
        FFS_RLOS_LO2    : out    vl_logic;
        FFS_RLOS_LO3    : out    vl_logic;
        ADDRI_7         : in     vl_logic;
        ADDRI_6         : in     vl_logic;
        ADDRI_5         : in     vl_logic;
        ADDRI_4         : in     vl_logic;
        ADDRI_3         : in     vl_logic;
        ADDRI_2         : in     vl_logic;
        ADDRI_1         : in     vl_logic;
        ADDRI_0         : in     vl_logic;
        WDATAI_7        : in     vl_logic;
        WDATAI_6        : in     vl_logic;
        WDATAI_5        : in     vl_logic;
        WDATAI_4        : in     vl_logic;
        WDATAI_3        : in     vl_logic;
        WDATAI_2        : in     vl_logic;
        WDATAI_1        : in     vl_logic;
        WDATAI_0        : in     vl_logic;
        RDI             : in     vl_logic;
        WSTBI           : in     vl_logic;
        CS_CHIF_0       : in     vl_logic;
        CS_CHIF_1       : in     vl_logic;
        CS_CHIF_2       : in     vl_logic;
        CS_CHIF_3       : in     vl_logic;
        CS_QIF          : in     vl_logic;
        QUAD_ID_1       : in     vl_logic;
        QUAD_ID_0       : in     vl_logic;
        RDATAO_7        : out    vl_logic;
        RDATAO_6        : out    vl_logic;
        RDATAO_5        : out    vl_logic;
        RDATAO_4        : out    vl_logic;
        RDATAO_3        : out    vl_logic;
        RDATAO_2        : out    vl_logic;
        RDATAO_1        : out    vl_logic;
        RDATAO_0        : out    vl_logic;
        INTO            : out    vl_logic;
        FF_SYSCLK_P1    : out    vl_logic;
        FF_SYSCLK0      : out    vl_logic;
        FF_SYSCLK1      : out    vl_logic;
        FF_SYSCLK2      : out    vl_logic;
        FF_SYSCLK3      : out    vl_logic;
        FF_RXCLK_P1     : out    vl_logic;
        FF_RXCLK_P2     : out    vl_logic;
        FF_RXCLK0       : out    vl_logic;
        FF_RXCLK1       : out    vl_logic;
        FF_RXCLK2       : out    vl_logic;
        FF_RXCLK3       : out    vl_logic;
        QUAD_CLK        : out    vl_logic;
        GRP_CLK_P1_3    : in     vl_logic;
        GRP_CLK_P1_2    : in     vl_logic;
        GRP_CLK_P1_1    : in     vl_logic;
        GRP_CLK_P1_0    : in     vl_logic;
        GRP_CLK_P2_3    : in     vl_logic;
        GRP_CLK_P2_2    : in     vl_logic;
        GRP_CLK_P2_1    : in     vl_logic;
        GRP_CLK_P2_0    : in     vl_logic;
        GRP_START_3     : in     vl_logic;
        GRP_START_2     : in     vl_logic;
        GRP_START_1     : in     vl_logic;
        GRP_START_0     : in     vl_logic;
        GRP_DONE_3      : in     vl_logic;
        GRP_DONE_2      : in     vl_logic;
        GRP_DONE_1      : in     vl_logic;
        GRP_DONE_0      : in     vl_logic;
        GRP_DESKEW_ERROR_3: in     vl_logic;
        GRP_DESKEW_ERROR_2: in     vl_logic;
        GRP_DESKEW_ERROR_1: in     vl_logic;
        GRP_DESKEW_ERROR_0: in     vl_logic;
        IQA_START_LS    : out    vl_logic;
        IQA_DONE_LS     : out    vl_logic;
        IQA_AND_FP1_LS  : out    vl_logic;
        IQA_AND_FP0_LS  : out    vl_logic;
        IQA_OR_FP1_LS   : out    vl_logic;
        IQA_OR_FP0_LS   : out    vl_logic;
        IQA_RST_N       : out    vl_logic;
        FFC_CK_CORE_TX  : in     vl_logic;
        FFC_CK_CORE_RX  : in     vl_logic;
        FF_TCLK0        : in     vl_logic;
        FF_TCLK1        : in     vl_logic;
        FF_TCLK2        : in     vl_logic;
        FF_TCLK3        : in     vl_logic;
        FF_RCLK0        : in     vl_logic;
        FF_RCLK1        : in     vl_logic;
        FF_RCLK2        : in     vl_logic;
        FF_RCLK3        : in     vl_logic;
        FF_TXD_0_23     : in     vl_logic;
        FF_TXD_0_22     : in     vl_logic;
        FF_TXD_0_21     : in     vl_logic;
        FF_TXD_0_20     : in     vl_logic;
        FF_TXD_0_19     : in     vl_logic;
        FF_TXD_0_18     : in     vl_logic;
        FF_TXD_0_17     : in     vl_logic;
        FF_TXD_0_16     : in     vl_logic;
        FF_TXD_0_15     : in     vl_logic;
        FF_TXD_0_14     : in     vl_logic;
        FF_TXD_0_13     : in     vl_logic;
        FF_TXD_0_12     : in     vl_logic;
        FF_TXD_0_11     : in     vl_logic;
        FF_TXD_0_10     : in     vl_logic;
        FF_TXD_0_9      : in     vl_logic;
        FF_TXD_0_8      : in     vl_logic;
        FF_TXD_0_7      : in     vl_logic;
        FF_TXD_0_6      : in     vl_logic;
        FF_TXD_0_5      : in     vl_logic;
        FF_TXD_0_4      : in     vl_logic;
        FF_TXD_0_3      : in     vl_logic;
        FF_TXD_0_2      : in     vl_logic;
        FF_TXD_0_1      : in     vl_logic;
        FF_TXD_0_0      : in     vl_logic;
        FF_TXD_1_23     : in     vl_logic;
        FF_TXD_1_22     : in     vl_logic;
        FF_TXD_1_21     : in     vl_logic;
        FF_TXD_1_20     : in     vl_logic;
        FF_TXD_1_19     : in     vl_logic;
        FF_TXD_1_18     : in     vl_logic;
        FF_TXD_1_17     : in     vl_logic;
        FF_TXD_1_16     : in     vl_logic;
        FF_TXD_1_15     : in     vl_logic;
        FF_TXD_1_14     : in     vl_logic;
        FF_TXD_1_13     : in     vl_logic;
        FF_TXD_1_12     : in     vl_logic;
        FF_TXD_1_11     : in     vl_logic;
        FF_TXD_1_10     : in     vl_logic;
        FF_TXD_1_9      : in     vl_logic;
        FF_TXD_1_8      : in     vl_logic;
        FF_TXD_1_7      : in     vl_logic;
        FF_TXD_1_6      : in     vl_logic;
        FF_TXD_1_5      : in     vl_logic;
        FF_TXD_1_4      : in     vl_logic;
        FF_TXD_1_3      : in     vl_logic;
        FF_TXD_1_2      : in     vl_logic;
        FF_TXD_1_1      : in     vl_logic;
        FF_TXD_1_0      : in     vl_logic;
        FF_TXD_2_23     : in     vl_logic;
        FF_TXD_2_22     : in     vl_logic;
        FF_TXD_2_21     : in     vl_logic;
        FF_TXD_2_20     : in     vl_logic;
        FF_TXD_2_19     : in     vl_logic;
        FF_TXD_2_18     : in     vl_logic;
        FF_TXD_2_17     : in     vl_logic;
        FF_TXD_2_16     : in     vl_logic;
        FF_TXD_2_15     : in     vl_logic;
        FF_TXD_2_14     : in     vl_logic;
        FF_TXD_2_13     : in     vl_logic;
        FF_TXD_2_12     : in     vl_logic;
        FF_TXD_2_11     : in     vl_logic;
        FF_TXD_2_10     : in     vl_logic;
        FF_TXD_2_9      : in     vl_logic;
        FF_TXD_2_8      : in     vl_logic;
        FF_TXD_2_7      : in     vl_logic;
        FF_TXD_2_6      : in     vl_logic;
        FF_TXD_2_5      : in     vl_logic;
        FF_TXD_2_4      : in     vl_logic;
        FF_TXD_2_3      : in     vl_logic;
        FF_TXD_2_2      : in     vl_logic;
        FF_TXD_2_1      : in     vl_logic;
        FF_TXD_2_0      : in     vl_logic;
        FF_TXD_3_23     : in     vl_logic;
        FF_TXD_3_22     : in     vl_logic;
        FF_TXD_3_21     : in     vl_logic;
        FF_TXD_3_20     : in     vl_logic;
        FF_TXD_3_19     : in     vl_logic;
        FF_TXD_3_18     : in     vl_logic;
        FF_TXD_3_17     : in     vl_logic;
        FF_TXD_3_16     : in     vl_logic;
        FF_TXD_3_15     : in     vl_logic;
        FF_TXD_3_14     : in     vl_logic;
        FF_TXD_3_13     : in     vl_logic;
        FF_TXD_3_12     : in     vl_logic;
        FF_TXD_3_11     : in     vl_logic;
        FF_TXD_3_10     : in     vl_logic;
        FF_TXD_3_9      : in     vl_logic;
        FF_TXD_3_8      : in     vl_logic;
        FF_TXD_3_7      : in     vl_logic;
        FF_TXD_3_6      : in     vl_logic;
        FF_TXD_3_5      : in     vl_logic;
        FF_TXD_3_4      : in     vl_logic;
        FF_TXD_3_3      : in     vl_logic;
        FF_TXD_3_2      : in     vl_logic;
        FF_TXD_3_1      : in     vl_logic;
        FF_TXD_3_0      : in     vl_logic;
        TCK_FMACP       : in     vl_logic;
        TESTCLK_MACO    : in     vl_logic;
        FB_RXD_0_23     : out    vl_logic;
        FB_RXD_0_22     : out    vl_logic;
        FB_RXD_0_21     : out    vl_logic;
        FB_RXD_0_20     : out    vl_logic;
        FB_RXD_0_19     : out    vl_logic;
        FB_RXD_0_18     : out    vl_logic;
        FB_RXD_0_17     : out    vl_logic;
        FB_RXD_0_16     : out    vl_logic;
        FB_RXD_0_15     : out    vl_logic;
        FB_RXD_0_14     : out    vl_logic;
        FB_RXD_0_13     : out    vl_logic;
        FB_RXD_0_12     : out    vl_logic;
        FB_RXD_0_11     : out    vl_logic;
        FB_RXD_0_10     : out    vl_logic;
        FB_RXD_0_9      : out    vl_logic;
        FB_RXD_0_8      : out    vl_logic;
        FB_RXD_0_7      : out    vl_logic;
        FB_RXD_0_6      : out    vl_logic;
        FB_RXD_0_5      : out    vl_logic;
        FB_RXD_0_4      : out    vl_logic;
        FB_RXD_0_3      : out    vl_logic;
        FB_RXD_0_2      : out    vl_logic;
        FB_RXD_0_1      : out    vl_logic;
        FB_RXD_0_0      : out    vl_logic;
        FB_RXD_1_23     : out    vl_logic;
        FB_RXD_1_22     : out    vl_logic;
        FB_RXD_1_21     : out    vl_logic;
        FB_RXD_1_20     : out    vl_logic;
        FB_RXD_1_19     : out    vl_logic;
        FB_RXD_1_18     : out    vl_logic;
        FB_RXD_1_17     : out    vl_logic;
        FB_RXD_1_16     : out    vl_logic;
        FB_RXD_1_15     : out    vl_logic;
        FB_RXD_1_14     : out    vl_logic;
        FB_RXD_1_13     : out    vl_logic;
        FB_RXD_1_12     : out    vl_logic;
        FB_RXD_1_11     : out    vl_logic;
        FB_RXD_1_10     : out    vl_logic;
        FB_RXD_1_9      : out    vl_logic;
        FB_RXD_1_8      : out    vl_logic;
        FB_RXD_1_7      : out    vl_logic;
        FB_RXD_1_6      : out    vl_logic;
        FB_RXD_1_5      : out    vl_logic;
        FB_RXD_1_4      : out    vl_logic;
        FB_RXD_1_3      : out    vl_logic;
        FB_RXD_1_2      : out    vl_logic;
        FB_RXD_1_1      : out    vl_logic;
        FB_RXD_1_0      : out    vl_logic;
        FB_RXD_2_23     : out    vl_logic;
        FB_RXD_2_22     : out    vl_logic;
        FB_RXD_2_21     : out    vl_logic;
        FB_RXD_2_20     : out    vl_logic;
        FB_RXD_2_19     : out    vl_logic;
        FB_RXD_2_18     : out    vl_logic;
        FB_RXD_2_17     : out    vl_logic;
        FB_RXD_2_16     : out    vl_logic;
        FB_RXD_2_15     : out    vl_logic;
        FB_RXD_2_14     : out    vl_logic;
        FB_RXD_2_13     : out    vl_logic;
        FB_RXD_2_12     : out    vl_logic;
        FB_RXD_2_11     : out    vl_logic;
        FB_RXD_2_10     : out    vl_logic;
        FB_RXD_2_9      : out    vl_logic;
        FB_RXD_2_8      : out    vl_logic;
        FB_RXD_2_7      : out    vl_logic;
        FB_RXD_2_6      : out    vl_logic;
        FB_RXD_2_5      : out    vl_logic;
        FB_RXD_2_4      : out    vl_logic;
        FB_RXD_2_3      : out    vl_logic;
        FB_RXD_2_2      : out    vl_logic;
        FB_RXD_2_1      : out    vl_logic;
        FB_RXD_2_0      : out    vl_logic;
        FB_RXD_3_23     : out    vl_logic;
        FB_RXD_3_22     : out    vl_logic;
        FB_RXD_3_21     : out    vl_logic;
        FB_RXD_3_20     : out    vl_logic;
        FB_RXD_3_19     : out    vl_logic;
        FB_RXD_3_18     : out    vl_logic;
        FB_RXD_3_17     : out    vl_logic;
        FB_RXD_3_16     : out    vl_logic;
        FB_RXD_3_15     : out    vl_logic;
        FB_RXD_3_14     : out    vl_logic;
        FB_RXD_3_13     : out    vl_logic;
        FB_RXD_3_12     : out    vl_logic;
        FB_RXD_3_11     : out    vl_logic;
        FB_RXD_3_10     : out    vl_logic;
        FB_RXD_3_9      : out    vl_logic;
        FB_RXD_3_8      : out    vl_logic;
        FB_RXD_3_7      : out    vl_logic;
        FB_RXD_3_6      : out    vl_logic;
        FB_RXD_3_5      : out    vl_logic;
        FB_RXD_3_4      : out    vl_logic;
        FB_RXD_3_3      : out    vl_logic;
        FB_RXD_3_2      : out    vl_logic;
        FB_RXD_3_1      : out    vl_logic;
        FB_RXD_3_0      : out    vl_logic;
        TCK_FMAC        : out    vl_logic;
        BS4PAD_0        : out    vl_logic;
        BS4PAD_1        : out    vl_logic;
        BS4PAD_2        : out    vl_logic;
        BS4PAD_3        : out    vl_logic;
        COUT_21         : out    vl_logic;
        COUT_20         : out    vl_logic;
        COUT_19         : out    vl_logic;
        COUT_18         : out    vl_logic;
        COUT_17         : out    vl_logic;
        COUT_16         : out    vl_logic;
        COUT_15         : out    vl_logic;
        COUT_14         : out    vl_logic;
        COUT_13         : out    vl_logic;
        COUT_12         : out    vl_logic;
        COUT_11         : out    vl_logic;
        COUT_10         : out    vl_logic;
        COUT_9          : out    vl_logic;
        COUT_8          : out    vl_logic;
        COUT_7          : out    vl_logic;
        COUT_6          : out    vl_logic;
        COUT_5          : out    vl_logic;
        COUT_4          : out    vl_logic;
        COUT_3          : out    vl_logic;
        COUT_2          : out    vl_logic;
        COUT_1          : out    vl_logic;
        COUT_0          : out    vl_logic;
        CIN_12          : in     vl_logic;
        CIN_11          : in     vl_logic;
        CIN_10          : in     vl_logic;
        CIN_9           : in     vl_logic;
        CIN_8           : in     vl_logic;
        CIN_7           : in     vl_logic;
        CIN_6           : in     vl_logic;
        CIN_5           : in     vl_logic;
        CIN_4           : in     vl_logic;
        CIN_3           : in     vl_logic;
        CIN_2           : in     vl_logic;
        CIN_1           : in     vl_logic;
        CIN_0           : in     vl_logic
    );
end PCSA_sim;
