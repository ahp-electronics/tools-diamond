library verilog;
use verilog.vl_types.all;
entity config_core_clocks is
    port(
        scanen          : in     vl_logic;
        wb_clk_nt       : in     vl_logic;
        smclk_tree      : out    vl_logic;
        smclk_tree_scan_off: out    vl_logic;
        hse_clk         : out    vl_logic;
        mx_smclk        : out    vl_logic;
        smclk_ext       : out    vl_logic;
        smclk_int       : out    vl_logic;
        smclk_div       : in     vl_logic;
        hse_clk_div     : in     vl_logic;
        sedclk          : out    vl_logic;
        cib_sed_clk     : in     vl_logic;
        sedclk_div      : in     vl_logic;
        sedclk_int_sel  : in     vl_logic;
        i2c_clk_prm     : out    vl_logic;
        isc_operational : in     vl_logic;
        fast_intclk     : out    vl_logic;
        slow_intclk     : out    vl_logic;
        intclk          : in     vl_logic;
        mclk_int        : out    vl_logic;
        mfg_tckmclk     : in     vl_logic;
        mclk_div        : in     vl_logic;
        mclk_byp        : out    vl_logic;
        mclk_byp_sel    : in     vl_logic_vector(1 downto 0);
        jtck            : out    vl_logic;
        mfg_clk_obsv_sel: in     vl_logic_vector(1 downto 0);
        tck_tree        : out    vl_logic;
        tck_pin         : in     vl_logic;
        rti_npd         : in     vl_logic;
        scpu_writen     : in     vl_logic;
        smclk_sel_enc   : in     vl_logic_vector(1 downto 0);
        jtag_disable    : in     vl_logic;
        sram_asr_clk    : out    vl_logic;
        dsr_clk         : out    vl_logic;
        tdr_sel_tck     : in     vl_logic;
        sck_tcv         : out    vl_logic;
        cclk_pin        : in     vl_logic;
        enable_cclk     : in     vl_logic;
        sspi_holdn      : in     vl_logic;
        njtrx_rst_async : in     vl_logic;
        persist_mspi    : in     vl_logic;
        mclk_pin        : in     vl_logic;
        mclk_en         : in     vl_logic;
        mclk_pol        : in     vl_logic;
        sck_tcv_sel     : in     vl_logic_vector(1 downto 0);
        scl_in_pad      : in     vl_logic;
        scl_clk_deb     : in     vl_logic;
        persist_i2c     : in     vl_logic;
        i2c_1st_addr_match_cfg: in     vl_logic;
        wbcact          : in     vl_logic;
        fifo_clk        : out    vl_logic;
        fifo_clk_sel    : in     vl_logic_vector(1 downto 0);
        i2c_2nd_scl_clk : out    vl_logic;
        scl_in_cib      : in     vl_logic;
        i2c_1st_scl_clk : out    vl_logic;
        spi_port_sck_tcv: out    vl_logic;
        spi_port_sck_tcv_inv: in     vl_logic;
        spi2nd_men      : in     vl_logic;
        sclk_i_2nd      : in     vl_logic;
        wkupclk         : out    vl_logic;
        cib_wkup_clk    : in     vl_logic;
        cib_wkup_clk_sel: in     vl_logic
    );
end config_core_clocks;
