library verilog;
use verilog.vl_types.all;
entity ao_22222222 is
    port(
        A               : in     vl_logic_vector(7 downto 0);
        EN              : in     vl_logic_vector(7 downto 0);
        Z               : out    vl_logic
    );
end ao_22222222;
