library verilog;
use verilog.vl_types.all;
entity cfg_cdu is
    port(
        sfdp_en         : in     vl_logic;
        njbse_sign_read : in     vl_logic;
        njbse_sign_cmd  : in     vl_logic;
        njbse_sign_cmd_read: in     vl_logic;
        sign_match      : out    vl_logic;
        preamblePass    : out    vl_logic;
        signatureCheckEvent: out    vl_logic;
        INT_SPI_CTRL    : in     vl_logic_vector(1 downto 0);
        scanen          : in     vl_logic;
        smclk           : in     vl_logic;
        smclk_int       : in     vl_logic;
        smclk_ext       : in     vl_logic;
        sedclk          : in     vl_logic;
        fifo_clk        : in     vl_logic;
        sck_tcv         : in     vl_logic;
        mclk_byp        : in     vl_logic;
        i2c_clk_prm     : in     vl_logic;
        mclk_int        : in     vl_logic;
        spi_port_sck_tcv: in     vl_logic;
        por             : in     vl_logic;
        slow_intclk     : in     vl_logic;
        fast_intclk     : in     vl_logic;
        nj_rst_async    : in     vl_logic;
        nj_rst_sync     : in     vl_logic;
        nji2c_rst_async : in     vl_logic;
        njtrx_rst_async : in     vl_logic;
        njtrx_rst_async0: in     vl_logic;
        isc_operational : in     vl_logic;
        isc_exec_b      : in     vl_logic;
        isc_exec_e      : in     vl_logic;
        isc_disable_exec: in     vl_logic;
        cfg_i2c_dat     : in     vl_logic_vector(15 downto 0);
        lsc_i2ci_crbr_wt_qual: in     vl_logic;
        lsc_i2ci_txdr_wt_qual: in     vl_logic;
        lsc_i2ci_rxdr_rd_qual: in     vl_logic;
        lsc_i2ci_sr_rd_qual: in     vl_logic;
        njvfy_rst_exec  : in     vl_logic;
        isc_done        : in     vl_logic;
        wkup_done       : in     vl_logic;
        cib_wkupclk_en  : in     vl_logic;
        ref_sys_slow    : in     vl_logic;
        sed_en          : in     vl_logic;
        restart_bse_en  : in     vl_logic;
        njboot_dat      : in     vl_logic_vector(7 downto 0);
        jtag_active_smsync_jb: in     vl_logic;
        tck_pin         : in     vl_logic;
        tck             : in     vl_logic;
        tdi             : in     vl_logic;
        cclk_in         : in     vl_logic;
        mclk_in         : in     vl_logic;
        scm_si          : in     vl_logic;
        sspi_si         : in     vl_logic;
        sspi_csn        : in     vl_logic;
        sspi_holdn      : in     vl_logic;
        scpu_csn        : in     vl_logic;
        scpu_writen     : in     vl_logic;
        din_16          : in     vl_logic_vector(15 downto 0);
        programn_pin    : in     vl_logic;
        initn_pin       : in     vl_logic;
        done_pin        : in     vl_logic;
        gsrn_pin        : in     vl_logic;
        cfg_pin         : in     vl_logic_vector(2 downto 0);
        mspisel_pin     : in     vl_logic_vector(3 downto 0);
        csn_pin         : in     vl_logic_vector(1 downto 0);
        sda_in_cfg      : in     vl_logic;
        scl_in_cfg      : in     vl_logic;
        sda_in_cib      : in     vl_logic;
        scl_in_cib      : in     vl_logic;
        sclk_i_2nd      : in     vl_logic;
        mosi_i_2nd      : in     vl_logic;
        miso_i_2nd      : in     vl_logic;
        scsn_2nd_cib    : in     vl_logic;
        rti             : in     vl_logic;
        seldr_ss        : in     vl_logic;
        shiftdr_ss      : in     vl_logic;
        updr_ss         : in     vl_logic;
        upir_ss         : in     vl_logic;
        exit1dr_ss      : in     vl_logic;
        ShiftDR         : in     vl_logic;
        tdrclk_sw_i     : in     vl_logic;
        busy_seldr      : in     vl_logic;
        jburst_en       : in     vl_logic;
        jburst_pause    : in     vl_logic;
        jburst_01       : in     vl_logic;
        jburst_08       : in     vl_logic;
        jpspi_en_norm   : in     vl_logic;
        jpspi_en_stack  : in     vl_logic;
        jpspi_en_int    : in     vl_logic;
        jpspi_param     : in     vl_logic_vector(7 downto 0);
        njshf_dat0      : in     vl_logic;
        njshf_dat_nd    : in     vl_logic;
        nj_rcv_rd_cmd   : in     vl_logic;
        njs_halt        : in     vl_logic;
        rfifo_re        : in     vl_logic;
        wfifo_we        : in     vl_logic;
        wfifo_din       : in     vl_logic_vector(7 downto 0);
        njpspi_en_norm  : in     vl_logic;
        njpspi_en_stack : in     vl_logic;
        njpspi_en_int   : in     vl_logic;
        njpspi_param    : in     vl_logic_vector(7 downto 0);
        ref_boot0       : in     vl_logic;
        ref_boot1       : in     vl_logic;
        ref_boot2       : in     vl_logic;
        initn_tmr       : in     vl_logic;
        goe_tmr         : in     vl_logic;
        done_tmr        : in     vl_logic;
        cfg_mstr_start  : in     vl_logic;
        cfg_mstr_stop   : in     vl_logic;
        njbse_sstcmd    : in     vl_logic;
        njbse_txcmd     : in     vl_logic;
        njbse_preamble  : in     vl_logic;
        njbse_rxall     : in     vl_logic;
        njbse_bypass    : in     vl_logic;
        njbse_fthrough  : in     vl_logic;
        tx_setmcpu      : in     vl_logic;
        tx_command      : in     vl_logic;
        tx_operand      : in     vl_logic;
        cfg_mtx_dat     : in     vl_logic_vector(7 downto 0);
        cfg_mcsn_dat    : in     vl_logic_vector(7 downto 0);
        ctrl_sspi_auto  : in     vl_logic;
        ctrl_cpu_manu   : in     vl_logic;
        ctrl_smfreq_sel : in     vl_logic_vector(1 downto 0);
        ctrl_hsefreq_sel: in     vl_logic_vector(1 downto 0);
        ctrl_hsediv2freq_sel: in     vl_logic;
        ctrl_mfreq_div  : in     vl_logic_vector(5 downto 0);
        ctrl_cpol       : in     vl_logic;
        ctrl_cpha       : in     vl_logic;
        ctrl_lsbf       : in     vl_logic;
        ctrl_mclk_byp   : in     vl_logic;
        ctrl_tx_edge    : in     vl_logic;
        ctrl_done_opt   : in     vl_logic_vector(1 downto 0);
        ctrl_initn_opt  : in     vl_logic_vector(1 downto 0);
        cfg_ctrl0_upd   : in     vl_logic;
        trim_sda_del    : in     vl_logic_vector(3 downto 0);
        pwr_save_mode   : in     vl_logic;
        mc1_dts_clk     : in     vl_logic;
        mc1_sync_source : in     vl_logic;
        mc1_sed_clk     : in     vl_logic_vector(6 downto 0);
        mc1_usr_clk     : in     vl_logic_vector(6 downto 0);
        cib_wkup_clk    : in     vl_logic;
        mfg_clkx2       : in     vl_logic;
        mfg_tckrti      : in     vl_logic;
        mfg_tckrti_force: in     vl_logic;
        mfg_tckmclk     : in     vl_logic;
        mfg_scpu_en     : in     vl_logic;
        int_spi_din     : in     vl_logic_vector(15 downto 0);
        sd_i2c_addr     : in     vl_logic_vector(7 downto 0);
        mc1_persist_mspi: in     vl_logic;
        mc1_persist_sspi: in     vl_logic;
        mc1_persist_i2c : in     vl_logic;
        mc1_persist_cpu8: in     vl_logic;
        mc1_persist_cpu16: in     vl_logic;
        fsd_persistn_progn: in     vl_logic;
        fsd_persist_initn: in     vl_logic;
        fsd_persist_done: in     vl_logic;
        fsd_persistn_sspi: in     vl_logic;
        fsd_persistn_i2c: in     vl_logic;
        fsd_persist_mspi: in     vl_logic;
        fsd_boot_sel    : in     vl_logic_vector(2 downto 0);
        mc1_persist_cap : in     vl_logic;
        cib_persist_in  : in     vl_logic_vector(15 downto 0);
        wb_clk_i        : in     vl_logic;
        spicr0          : in     vl_logic_vector(7 downto 0);
        spicr1          : in     vl_logic_vector(7 downto 0);
        spicr2          : in     vl_logic_vector(7 downto 0);
        spibr           : in     vl_logic_vector(7 downto 0);
        spicsr          : in     vl_logic_vector(7 downto 0);
        spitxdr         : in     vl_logic_vector(7 downto 0);
        wb_spicr0_wt    : in     vl_logic;
        wb_spicr1_wt    : in     vl_logic;
        wb_spicr2_wt    : in     vl_logic;
        wb_spibr_wt     : in     vl_logic;
        wb_spicsr_wt    : in     vl_logic;
        wb_spitxdr_wt   : in     vl_logic;
        wb_spirxdr_rd   : in     vl_logic;
        wbccr1          : in     vl_logic_vector(7 downto 0);
        wbctxdr         : in     vl_logic_vector(7 downto 0);
        wb_wbccr1_wt    : in     vl_logic;
        wb_wbctxdr_wt   : in     vl_logic;
        wb_wbcrxdr_rd   : in     vl_logic;
        i2ccr1_1st      : in     vl_logic_vector(7 downto 0);
        i2ccmdr_1st     : in     vl_logic_vector(7 downto 0);
        i2ctxdr_1st     : in     vl_logic_vector(7 downto 0);
        i2cbr_1st       : in     vl_logic_vector(9 downto 0);
        wb_i2ccr1_wt_1st: in     vl_logic;
        wb_i2ccmdr_wt_1st: in     vl_logic;
        wb_i2cbr_wt_1st : in     vl_logic;
        wb_i2ctxdr_wt_1st: in     vl_logic;
        wb_i2crxdr_rd_1st: in     vl_logic;
        wb_i2cgcdr_rd_1st: in     vl_logic;
        i2ccr1_2nd      : in     vl_logic_vector(7 downto 0);
        i2ccmdr_2nd     : in     vl_logic_vector(7 downto 0);
        i2ctxdr_2nd     : in     vl_logic_vector(7 downto 0);
        i2cbr_2nd       : in     vl_logic_vector(9 downto 0);
        wb_i2ccr1_wt_2nd: in     vl_logic;
        wb_i2ccmdr_wt_2nd: in     vl_logic;
        wb_i2cbr_wt_2nd : in     vl_logic;
        wb_i2ctxdr_wt_2nd: in     vl_logic;
        wb_i2crxdr_rd_2nd: in     vl_logic;
        wb_i2cgcdr_rd_2nd: in     vl_logic;
        cfg0_latter     : in     vl_logic;
        mcsn_o_1st      : out    vl_logic_vector(7 downto 0);
        mcsn_oe_1st     : out    vl_logic_vector(7 downto 0);
        mclk_o_1st      : out    vl_logic;
        mclk_oe_1st     : out    vl_logic;
        sspi_so_1st     : out    vl_logic;
        sspi_oe_1st     : out    vl_logic;
        mclk_byp_o      : out    vl_logic;
        mclk_byp_oe     : out    vl_logic;
        data_o_1st      : out    vl_logic_vector(15 downto 0);
        data_oe_1st     : out    vl_logic_vector(15 downto 0);
        docson_o        : out    vl_logic;
        docson_oe       : out    vl_logic;
        busy_o_1st      : out    vl_logic;
        busy_oe_1st     : out    vl_logic;
        initn_o         : out    vl_logic;
        initn_oe        : out    vl_logic;
        donep_o         : out    vl_logic;
        donep_oe        : out    vl_logic;
        persist_mspi    : out    vl_logic;
        persist_sspi    : out    vl_logic;
        persist_i2c     : out    vl_logic;
        persist_cpu8    : out    vl_logic;
        persist_cpu16   : out    vl_logic;
        p_slave         : out    vl_logic;
        p_scm           : out    vl_logic;
        p_scpu          : out    vl_logic;
        p_mspi0         : out    vl_logic;
        p_mspim         : out    vl_logic;
        p_mp8           : out    vl_logic;
        p_mp16          : out    vl_logic;
        p_mspi_slow     : out    vl_logic;
        p_mspi_fast     : out    vl_logic;
        p_mspi_dual     : out    vl_logic;
        p_mspi_quad     : out    vl_logic;
        p_mp8_quad      : out    vl_logic;
        p_mp16_quad     : out    vl_logic;
        p_mspi_all      : out    vl_logic;
        p_sst           : out    vl_logic;
        p_end_bpft      : out    vl_logic;
        p_eboot0p       : out    vl_logic;
        p_eboot1p       : out    vl_logic;
        p_eboot1s       : out    vl_logic;
        p_eboot2p       : out    vl_logic;
        p_eboot2s       : out    vl_logic;
        p_nboot         : out    vl_logic;
        p_iboot0p       : out    vl_logic;
        p_iboot1p       : out    vl_logic;
        p_iboot1s       : out    vl_logic;
        p_iboot2p       : out    vl_logic;
        p_iboot2s       : out    vl_logic;
        wbc_active      : out    vl_logic;
        sspi_active     : out    vl_logic;
        i2c_active      : out    vl_logic;
        extspi_out      : out    vl_logic;
        rfifo_out       : out    vl_logic_vector(7 downto 0);
        rfifo_empty     : out    vl_logic;
        rfifo_full      : out    vl_logic;
        rfifo_overflow  : out    vl_logic;
        wfifo_full      : out    vl_logic;
        wfifo_overflow  : out    vl_logic;
        cfg_mstr_busy   : out    vl_logic;
        njm_tr_next     : out    vl_logic;
        njm_tr_done     : out    vl_logic;
        njm_mcpu_done   : out    vl_logic;
        preamble_std    : out    vl_logic;
        preamble_enc    : out    vl_logic;
        preamble_std_ext: out    vl_logic;
        preamble_enc_ext: out    vl_logic;
        boot_setup      : out    vl_logic_vector(5 downto 0);
        cfg_i2c_dout    : out    vl_logic_vector(7 downto 0);
        programn_tog    : out    vl_logic;
        programn_pin_sync: out    vl_logic;
        initn_pin_sync  : out    vl_logic;
        done_pin_sync   : out    vl_logic;
        done_rise1      : out    vl_logic;
        gsrn_pin_sync   : out    vl_logic;
        njport_init     : out    vl_logic;
        njport_active   : out    vl_logic;
        njport_exec     : out    vl_logic;
        dtsclk          : out    vl_logic;
        usrclk          : out    vl_logic;
        int_spi_mclk    : out    vl_logic;
        int_spi_data    : out    vl_logic_vector(15 downto 0);
        int_spi_mcsn    : out    vl_logic_vector(7 downto 0);
        persist_out_cib : out    vl_logic_vector(15 downto 0);
        i2crxdr_1st     : out    vl_logic_vector(7 downto 0);
        i2cgcdr_1st     : out    vl_logic_vector(7 downto 0);
        i2csr_1st       : out    vl_logic_vector(7 downto 0);
        i2c_wkup_1st    : out    vl_logic;
        i2crxdr_2nd     : out    vl_logic_vector(7 downto 0);
        i2cgcdr_2nd     : out    vl_logic_vector(7 downto 0);
        i2csr_2nd       : out    vl_logic_vector(7 downto 0);
        i2c_wkup_2nd    : out    vl_logic;
        wbcsr           : out    vl_logic_vector(7 downto 0);
        wbcrxdr         : out    vl_logic_vector(7 downto 0);
        spisr           : out    vl_logic_vector(7 downto 0);
        spirxdr         : out    vl_logic_vector(7 downto 0);
        spi_wkup        : out    vl_logic;
        sda_out_cib     : out    vl_logic;
        sda_oe_cib      : out    vl_logic;
        scl_out_cib     : out    vl_logic;
        scl_oe_cib      : out    vl_logic;
        mcsn_o_cib      : out    vl_logic_vector(7 downto 0);
        mcsn_oe_cib     : out    vl_logic_vector(7 downto 0);
        mclk_o_2nd      : out    vl_logic;
        mclk_oe_2nd     : out    vl_logic;
        mosi_o_2nd      : out    vl_logic;
        mosi_oe_2nd     : out    vl_logic;
        miso_o_2nd      : out    vl_logic;
        miso_oe_2nd     : out    vl_logic;
        scl_clk_deb     : out    vl_logic;
        sda_out_cfg     : out    vl_logic;
        sda_oe_cfg      : out    vl_logic;
        scl_out_cfg     : out    vl_logic;
        scl_oe_cfg      : out    vl_logic;
        cfgmode_cfg     : out    vl_logic;
        cib_wkup_clk_sel: out    vl_logic;
        smclk_div       : out    vl_logic;
        hse_clk_div     : out    vl_logic;
        smclk_sel_enc   : out    vl_logic_vector(1 downto 0);
        rti_npd         : out    vl_logic;
        tdr_sel_tck     : out    vl_logic;
        sedclk_div      : out    vl_logic;
        mclk_div        : out    vl_logic;
        mclk_byp_sel    : out    vl_logic_vector(1 downto 0);
        sck_tcv_sel     : out    vl_logic_vector(1 downto 0);
        fifo_clk_sel    : out    vl_logic_vector(1 downto 0);
        wbcact          : out    vl_logic;
        mclk_en         : out    vl_logic;
        mclk_pol        : out    vl_logic;
        i2c_1st_addr_match_cfg: out    vl_logic;
        spi2nd_men      : out    vl_logic;
        spi_port_sck_tcv_inv: out    vl_logic;
        p_iboot0s       : out    vl_logic
    );
end cfg_cdu;
