library verilog;
use verilog.vl_types.all;
entity sbnx4v1mce_1 is
    port(
        A               : in     vl_logic;
        Z               : out    vl_logic
    );
end sbnx4v1mce_1;
