library verilog;
use verilog.vl_types.all;
entity vhim4mce is
    port(
        Z               : out    vl_logic
    );
end vhim4mce;
