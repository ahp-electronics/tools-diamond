library verilog;
use verilog.vl_types.all;
entity BOXT is
    port(
        USER_IRQ_OUT    : out    vl_logic;
        UPDTBSR         : out    vl_logic;
        TRI_ION         : out    vl_logic;
        TRESET          : out    vl_logic;
        TDOEN           : out    vl_logic;
        TDOE            : out    vl_logic;
        TDO             : out    vl_logic;
        TDI1_RASB       : out    vl_logic;
        TDI1_LASB       : out    vl_logic;
        TCK2            : out    vl_logic;
        SRI_WR          : out    vl_logic;
        SRI_WDATA       : out    vl_logic;
        SRI_RD          : out    vl_logic;
        SRI_CLK         : out    vl_logic;
        SRI_ADDR        : out    vl_logic_vector(9 downto 0);
        SPI_TRI_ION     : out    vl_logic;
        SHIFT_ADDR_2ND  : out    vl_logic;
        SHIFT_ADDR_1ST  : out    vl_logic;
        SHBSRN          : out    vl_logic;
        SERIAL_DATA     : out    vl_logic;
        RST_DATA_REG_N  : out    vl_logic;
        RST_ADDR_REG    : out    vl_logic;
        RDY_BUSY_N      : out    vl_logic;
        QOUT            : out    vl_logic;
        PWRUPRES        : out    vl_logic;
        PSRSFTN         : out    vl_logic;
        PSRENABLE3      : out    vl_logic;
        PSRENABLE2      : out    vl_logic;
        PSRENABLE1      : out    vl_logic;
        PSRCAP          : out    vl_logic;
        PRDY_TS         : out    vl_logic;
        PD7_3_TS        : out    vl_logic;
        PD31_16_TS      : out    vl_logic;
        PD2_0_TS        : out    vl_logic;
        PD15_8_TS       : out    vl_logic;
        PCS_SL_STRAIT   : out    vl_logic;
        PA_OUT          : out    vl_logic_vector(21 downto 0);
        MPI_TRI_ION     : out    vl_logic_vector(2 downto 0);
        MPI_DP_TS       : out    vl_logic_vector(2 downto 0);
        MPI_DP_TRI_ION  : out    vl_logic_vector(2 downto 0);
        MPI_CNTL_TS     : out    vl_logic;
        MPC_TEA         : out    vl_logic;
        MPC_TA          : out    vl_logic;
        MPC_RETRY       : out    vl_logic;
        MPC_RD_PARITY   : out    vl_logic_vector(0 to 3);
        LD_RDBKD        : out    vl_logic;
        LDC_N           : out    vl_logic;
        JUPDATE         : out    vl_logic;
        JTDI            : out    vl_logic;
        JSHIFT          : out    vl_logic;
        JRTI            : out    vl_logic_vector(8 downto 1);
        JRSTN           : out    vl_logic;
        JCE             : out    vl_logic_vector(8 downto 1);
        INTEST          : out    vl_logic;
        INIT_N          : out    vl_logic;
        INIT_1_DATA     : out    vl_logic;
        HSEL_RASBS      : out    vl_logic;
        HSEL_LASBS      : out    vl_logic;
        HIGHZ           : out    vl_logic;
        HDC             : out    vl_logic;
        HCLK_RASB       : out    vl_logic;
        HCLK_LASB       : out    vl_logic;
        HCLK_CIB        : out    vl_logic;
        GSR_N           : out    vl_logic;
        GSRN_SYNC       : out    vl_logic;
        GOT_DATA        : out    vl_logic;
        GOT_ADDR        : out    vl_logic;
        FSWRN           : out    vl_logic;
        FSWDATA         : out    vl_logic_vector(35 downto 0);
        FSSIZE          : out    vl_logic_vector(1 downto 0);
        FSRDY           : out    vl_logic;
        FSADDR          : out    vl_logic_vector(17 downto 0);
        FMRETRY         : out    vl_logic;
        FMRDATA         : out    vl_logic_vector(35 downto 0);
        FMERR           : out    vl_logic;
        FMACK           : out    vl_logic;
        EN_PDWN         : out    vl_logic;
        EN_OSC          : out    vl_logic;
        EN_CCLK_N       : out    vl_logic;
        EN_ADDR_INCR    : out    vl_logic;
        EN_ADDR         : out    vl_logic;
        ENTCK_JTAG      : out    vl_logic;
        DOUT            : out    vl_logic;
        DOBIST_RASB     : out    vl_logic;
        DOBIST_LASB     : out    vl_logic;
        DEBUG_BUS       : out    vl_logic_vector(15 downto 0);
        CPTBSR          : out    vl_logic;
        CFG_DATA_WR     : out    vl_logic;
        CFG_DATA_PC     : out    vl_logic;
        CFG_DATA        : out    vl_logic_vector(7 downto 0);
        CCLK_OUT        : out    vl_logic;
        CCLK_AD         : out    vl_logic;
        CAPTURE         : out    vl_logic;
        ADDR_TS         : out    vl_logic;
        MPC_RD_DATA     : out    vl_logic_vector(0 to 31);
        PAD_DONE        : out    vl_logic;
        CFG_CK          : out    vl_logic;
        PWR_ON          : out    vl_logic;
        DONE            : out    vl_logic;
        RDBK_DATA       : out    vl_logic;
        SRI_RST_N       : out    vl_logic;
        LASB_INIT_N     : out    vl_logic;
        RASB_INIT_N     : out    vl_logic;
        LASB_PWRUPRES   : out    vl_logic;
        RASB_PWRUPRES   : out    vl_logic;
        LASB_TRI_ION    : out    vl_logic;
        RASB_TRI_ION    : out    vl_logic;
        LASB_GSR_N      : out    vl_logic;
        RASB_GSR_N      : out    vl_logic;
        LASB_DONE       : out    vl_logic;
        RASB_DONE       : out    vl_logic;
        SYSB_DEBUG      : out    vl_logic_vector(23 downto 0);
        TCK_CIB         : out    vl_logic;
        TMS_CIB         : out    vl_logic;
        TDI_CIB         : out    vl_logic;
        BS_MODE         : out    vl_logic;
        SCANEN_LASB     : out    vl_logic;
        SCANEN_RASB     : out    vl_logic;
        TCK2_LASB       : out    vl_logic;
        TCK2_RASB       : out    vl_logic;
        TRESET_LASB     : out    vl_logic;
        TRESET_RASB     : out    vl_logic;
        PSRTRST         : out    vl_logic;
        SHDR_LASB       : out    vl_logic;
        SHDR_RASB       : out    vl_logic;
        CPTDR_LASB      : out    vl_logic;
        CPTDR_RASB      : out    vl_logic;
        RUNTST_LASB     : out    vl_logic;
        RUNTST_RASB     : out    vl_logic;
        UPDTDR_LASB     : out    vl_logic;
        UPDTDR_RASB     : out    vl_logic;
        JSCANENABLE     : out    vl_logic_vector(8 downto 1);
        JSCANIN         : out    vl_logic;
        TDI1            : out    vl_logic;
        JTCK            : out    vl_logic;
        J_BOXT_SCANEN   : out    vl_logic;
        SCANOUT         : out    vl_logic;
        BOXT_SE         : out    vl_logic;
        MPI_IRQ_N       : out    vl_logic;
        LASB_IRQ_OUT    : out    vl_logic;
        RASB_IRQ_OUT    : out    vl_logic;
        LASB_PAR_ODD    : out    vl_logic;
        RASB_PAR_ODD    : out    vl_logic;
        HRDATA_LASBM    : out    vl_logic_vector(35 downto 0);
        HRDATA_RASBM    : out    vl_logic_vector(35 downto 0);
        HWDATA_LASBS    : out    vl_logic_vector(35 downto 0);
        HWDATA_RASBS    : out    vl_logic_vector(35 downto 0);
        HADDR_LASBS     : out    vl_logic_vector(17 downto 0);
        HADDR_RASBS     : out    vl_logic_vector(17 downto 0);
        HTRANS_LASBS    : out    vl_logic_vector(1 downto 0);
        HTRANS_RASBS    : out    vl_logic_vector(1 downto 0);
        HRESP_LASBM     : out    vl_logic_vector(1 downto 0);
        HRESP_RASBM     : out    vl_logic_vector(1 downto 0);
        HSIZE_LASBS     : out    vl_logic_vector(1 downto 0);
        HSIZE_RASBS     : out    vl_logic_vector(1 downto 0);
        HBURST_LASBS    : out    vl_logic;
        HBURST_RASBS    : out    vl_logic;
        HRESET_N_LASB   : out    vl_logic;
        HRESET_N_RASB   : out    vl_logic;
        HGRANT_LASBM    : out    vl_logic;
        HGRANT_RASBM    : out    vl_logic;
        HWRITE_LASBS    : out    vl_logic;
        HWRITE_RASBS    : out    vl_logic;
        HREADY_LASB     : out    vl_logic;
        HREADY_RASB     : out    vl_logic;
        TIE_LOW         : out    vl_logic;
        TIE_HIGH        : out    vl_logic;
        BOXT_LOW        : out    vl_logic;
        BOXT_HIGH       : out    vl_logic;
        HCLK            : out    vl_logic;
        HRESET_N        : out    vl_logic;
        HREADY          : out    vl_logic;
        SBWR_O          : out    vl_logic_vector(33 downto 0);
        WR_N            : in     vl_logic;
        USR_TDO         : in     vl_logic;
        USR_START_CLK   : in     vl_logic;
        USR_GSR         : in     vl_logic;
        USR_CLK         : in     vl_logic;
        USER_IRQ_IN     : in     vl_logic;
        TS_ALL          : in     vl_logic;
        TMS             : in     vl_logic;
        TDI             : in     vl_logic;
        TCK             : in     vl_logic;
        SYS_RST_N       : in     vl_logic;
        SRI_RDATA       : in     vl_logic_vector(63 downto 0);
        SO_BIST_RASB    : in     vl_logic;
        SO_BIST_LASB    : in     vl_logic;
        SED_CLK         : in     vl_logic;
        RD_N            : in     vl_logic;
        RD_CFG_USR      : in     vl_logic;
        RD_CFG          : in     vl_logic;
        RDBK_ZERO_ALL_N : in     vl_logic;
        RDBK_DOUT       : in     vl_logic_vector(7 downto 0);
        RASB_SLAVE_ENABLE: in     vl_logic;
        RASB_SEL        : in     vl_logic;
        RASB_CLK        : in     vl_logic;
        PWRUP_NPUR      : in     vl_logic;
        PWRUP_E9        : in     vl_logic;
        PTEST_N         : in     vl_logic;
        PSROUT3         : in     vl_logic;
        PSROUT2         : in     vl_logic;
        PSROUT1         : in     vl_logic;
        MPI_RST_N       : in     vl_logic;
        MPI_CLK         : in     vl_logic;
        MPC_WR_PARITY   : in     vl_logic_vector(0 to 3);
        MPC_WR_DATA     : in     vl_logic_vector(0 to 31);
        MPC_TSIZ        : in     vl_logic_vector(0 to 1);
        MPC_BURST       : in     vl_logic;
        MPC_BDIP        : in     vl_logic;
        MPC_ADDR        : in     vl_logic_vector(14 to 31);
        MODE            : in     vl_logic_vector(3 downto 0);
        MC1_USR_TDO     : in     vl_logic;
        MC1_USR_SL      : in     vl_logic_vector(1 downto 0);
        MC1_USR_MR      : in     vl_logic_vector(1 downto 0);
        MC1_USR_CLK     : in     vl_logic;
        MC1_USERBIT     : in     vl_logic_vector(31 downto 0);
        MC1_USER        : in     vl_logic;
        MC1_TRI         : in     vl_logic_vector(3 downto 0);
        MC1_TIMEOUT_INDEX2: in     vl_logic_vector(3 downto 0);
        MC1_TIMEOUT_INDEX1: in     vl_logic_vector(3 downto 0);
        MC1_TEST_CTR    : in     vl_logic;
        MC1_SYS_RST     : in     vl_logic;
        MC1_STRT        : in     vl_logic_vector(4 downto 0);
        MC1_SPI_ADDR    : in     vl_logic_vector(31 downto 0);
        MC1_SED_CLK     : in     vl_logic;
        MC1_SCLK        : in     vl_logic;
        MC1_SCAN        : in     vl_logic_vector(8 downto 1);
        MC1_RST_RAM_N   : in     vl_logic;
        MC1_RST_HCLK_N  : in     vl_logic;
        MC1_RST_GSRN    : in     vl_logic;
        MC1_RST_BUS_N   : in     vl_logic;
        MC1_RDBK_REG    : in     vl_logic;
        MC1_PRIORITY_MPI: in     vl_logic_vector(1 downto 0);
        MC1_PRIORITY_FPGA: in     vl_logic_vector(1 downto 0);
        MC1_PRIORITY_ASB: in     vl_logic_vector(1 downto 0);
        MC1_PAR_ODD     : in     vl_logic;
        MC1_OSC_DIV     : in     vl_logic_vector(2 downto 0);
        MC1_OSC_CLK     : in     vl_logic;
        MC1_MPI_RST     : in     vl_logic;
        MC1_MPI_CLK     : in     vl_logic;
        MC1_MPI_ASYNC   : in     vl_logic;
        MC1_MPI         : in     vl_logic;
        MC1_MODE        : in     vl_logic_vector(3 downto 0);
        MC1_INTERRUPT_VECTOR_6: in     vl_logic_vector(31 downto 0);
        MC1_INTERRUPT_VECTOR_5: in     vl_logic_vector(31 downto 0);
        MC1_INTERRUPT_VECTOR_4: in     vl_logic_vector(31 downto 0);
        MC1_INTERRUPT_VECTOR_3: in     vl_logic_vector(31 downto 0);
        MC1_INTERRUPT_VECTOR_2: in     vl_logic_vector(31 downto 0);
        MC1_INTERRUPT_VECTOR_1: in     vl_logic_vector(31 downto 0);
        MC1_GSRN_SYNC   : in     vl_logic;
        MC1_GSRN_INV    : in     vl_logic;
        MC1_FPSC_CLK    : in     vl_logic;
        MC1_FPSC        : in     vl_logic;
        MC1_EXT_CCLK    : in     vl_logic;
        MC1_EN_SPI_N    : in     vl_logic;
        MC1_EN_SED      : in     vl_logic;
        MC1_EN_READCAP  : in     vl_logic;
        MC1_EN_RDBK     : in     vl_logic;
        MC1_EN_OSC      : in     vl_logic;
        MC1_EN_ONCE     : in     vl_logic;
        MC1_EN_MPI_PARITY: in     vl_logic;
        MC1_EN_CAPTURE  : in     vl_logic;
        MC1_DONE        : in     vl_logic_vector(1 downto 0);
        MC1_DIS_MODES   : in     vl_logic;
        LAST_ADDR       : in     vl_logic_vector(13 downto 0);
        LASB_SLAVE_ENABLE: in     vl_logic;
        LASB_CLK        : in     vl_logic;
        JTDO            : in     vl_logic_vector(8 downto 1);
        INITIN_N        : in     vl_logic;
        HRESP_RASBS     : in     vl_logic_vector(1 downto 0);
        HRESP_LASBS     : in     vl_logic_vector(1 downto 0);
        HREADY_RASBS    : in     vl_logic;
        HREADY_LASBS    : in     vl_logic;
        HRDATA_RASBS    : in     vl_logic_vector(35 downto 0);
        HRDATA_LASBS    : in     vl_logic_vector(35 downto 0);
        FSRETRY         : in     vl_logic;
        FSRESET_N       : in     vl_logic;
        FSRDATA         : in     vl_logic_vector(35 downto 0);
        FSIRQ           : in     vl_logic;
        FSERR           : in     vl_logic;
        FSCLK           : in     vl_logic;
        FSACK           : in     vl_logic;
        FMWRN           : in     vl_logic;
        FMWDATA         : in     vl_logic_vector(35 downto 0);
        FMSIZE          : in     vl_logic_vector(1 downto 0);
        FMRESET_N       : in     vl_logic;
        FMRDY           : in     vl_logic;
        FMLOCK          : in     vl_logic;
        FMIRQ           : in     vl_logic;
        FMCLK           : in     vl_logic;
        FMBURST         : in     vl_logic;
        FMADDR          : in     vl_logic_vector(17 downto 0);
        DONEIN          : in     vl_logic;
        DMA_TRI_DATA    : in     vl_logic;
        DMA_TRI_CTL     : in     vl_logic;
        DMA_TEA         : in     vl_logic;
        DMA_TA          : in     vl_logic;
        DMA_RETRY       : in     vl_logic;
        DMA_RD_PARITY   : in     vl_logic_vector(0 to 3);
        DMA_RD_DATA     : in     vl_logic_vector(0 to 31);
        CS1             : in     vl_logic;
        CS0_N           : in     vl_logic;
        CODE7           : in     vl_logic_vector(7 downto 0);
        CODE6           : in     vl_logic_vector(7 downto 0);
        CODE5           : in     vl_logic_vector(7 downto 0);
        CODE4           : in     vl_logic_vector(7 downto 0);
        CODE3           : in     vl_logic_vector(7 downto 0);
        CODE2           : in     vl_logic_vector(7 downto 0);
        CODE1           : in     vl_logic_vector(7 downto 0);
        CODE0           : in     vl_logic_vector(7 downto 0);
        CHIPID          : in     vl_logic_vector(7 downto 0);
        CFG_RESET_N     : in     vl_logic;
        CFG_PRGM_N      : in     vl_logic;
        CFG_OSC         : in     vl_logic;
        CCLKIN          : in     vl_logic;
        CAPT_I_N        : in     vl_logic;
        BSRSO           : in     vl_logic;
        ADDR_HIGH_DEL_N : in     vl_logic;
        PARTID          : in     vl_logic_vector(31 downto 0);
        SYS_SE          : in     vl_logic;
        BOXT_SFTEN      : in     vl_logic;
        SCANIN          : in     vl_logic;
        ENTCK           : in     vl_logic;
        SCANEN          : in     vl_logic;
        HWDATA_LASBM    : in     vl_logic_vector(35 downto 0);
        HWDATA_RASBM    : in     vl_logic_vector(35 downto 0);
        HADDR_LASBM     : in     vl_logic_vector(17 downto 0);
        HADDR_RASBM     : in     vl_logic_vector(17 downto 0);
        HTRANS_LASBM    : in     vl_logic_vector(1 downto 0);
        HTRANS_RASBM    : in     vl_logic_vector(1 downto 0);
        HSIZE_LASBM     : in     vl_logic_vector(1 downto 0);
        HSIZE_RASBM     : in     vl_logic_vector(1 downto 0);
        HBURST_LASBM    : in     vl_logic;
        HBURST_RASBM    : in     vl_logic;
        HBUSREQ_LASBM   : in     vl_logic;
        HBUSREQ_RASBM   : in     vl_logic;
        HLOCK_LASBM     : in     vl_logic;
        HLOCK_RASBM     : in     vl_logic;
        HWRITE_LASBM    : in     vl_logic;
        HWRITE_RASBM    : in     vl_logic;
        SCANOUT_LASB    : in     vl_logic;
        SCANOUT_RASB    : in     vl_logic;
        J_BOXT_SCANOUT  : in     vl_logic;
        LASB_IRQ_SLAVE  : in     vl_logic;
        RASB_IRQ_SLAVE  : in     vl_logic;
        LASB_IRQ_MASTER : in     vl_logic;
        RASB_IRQ_MASTER : in     vl_logic;
        LASB_GSR        : in     vl_logic;
        RASB_GSR        : in     vl_logic;
        TIELOW          : in     vl_logic;
        TIEHIGH         : in     vl_logic
    );
end BOXT;
