library verilog;
use verilog.vl_types.all;
entity MIPIDPHYA is
    generic(
        HSEL            : integer := 1;
        HS_16BIT_EN     : integer := 1;
        CN              : integer := 0;
        CM              : integer := 0;
        CO              : integer := 0;
        PLL_TST         : integer := 9;
        ENP_DESER       : integer := 0
    );
    port(
        CKP             : inout  vl_logic;
        CKN             : inout  vl_logic;
        CLKHSBYTE       : out    vl_logic;
        CLKRXHSEN       : in     vl_logic;
        CLKDRXLPP       : out    vl_logic;
        CLKRXLPEN       : in     vl_logic;
        CLKDRXLPN       : out    vl_logic;
        CLKCDEN         : in     vl_logic;
        CLKDCDN         : out    vl_logic;
        CLKDTXLPP       : in     vl_logic;
        CLKTXLPEN       : in     vl_logic;
        CLKDTXLPN       : in     vl_logic;
        CLKTXHSEN       : in     vl_logic;
        CLKTXHSGATE     : in     vl_logic;
        CLKTXHSPD       : in     vl_logic;
        CLKDRXHS        : out    vl_logic;
        HSBYTECLKD      : out    vl_logic;
        HSBYTECLKS      : out    vl_logic;
        LBEN            : in     vl_logic;
        PDDPHY          : in     vl_logic;
        PDBIAS          : in     vl_logic;
        PDCKG           : in     vl_logic;
        CLKREF          : in     vl_logic;
        LOCK            : out    vl_logic;
        PDPLL           : in     vl_logic;
        DP0             : inout  vl_logic;
        DP1             : inout  vl_logic;
        DP2             : inout  vl_logic;
        DP3             : inout  vl_logic;
        DN0             : inout  vl_logic;
        DN1             : inout  vl_logic;
        DN2             : inout  vl_logic;
        DN3             : inout  vl_logic;
        D0DRXLPP        : out    vl_logic;
        D0RXLPEN        : in     vl_logic;
        D0DRXLPN        : out    vl_logic;
        D0DCDP          : out    vl_logic;
        D0CDEN          : in     vl_logic;
        D0DCDN          : out    vl_logic;
        D0DTXLPP        : in     vl_logic;
        D0TXLPEN        : in     vl_logic;
        D0DTXLPN        : in     vl_logic;
        D0RXHSEN        : in     vl_logic;
        D0HSRXDATA15    : out    vl_logic;
        D0HSRXDATA14    : out    vl_logic;
        D0HSRXDATA13    : out    vl_logic;
        D0HSRXDATA12    : out    vl_logic;
        D0HSRXDATA11    : out    vl_logic;
        D0HSRXDATA10    : out    vl_logic;
        D0HSRXDATA9     : out    vl_logic;
        D0HSRXDATA8     : out    vl_logic;
        D0HSRXDATA7     : out    vl_logic;
        D0HSRXDATA6     : out    vl_logic;
        D0HSRXDATA5     : out    vl_logic;
        D0HSRXDATA4     : out    vl_logic;
        D0HSRXDATA3     : out    vl_logic;
        D0HSRXDATA2     : out    vl_logic;
        D0HSRXDATA1     : out    vl_logic;
        D0HSRXDATA0     : out    vl_logic;
        D0SYNC          : out    vl_logic;
        D0ERRSYNC       : out    vl_logic;
        D0NOSYNC        : out    vl_logic;
        D0HSDESEREN     : in     vl_logic;
        D0TXHSEN        : in     vl_logic;
        D0HSTXDATA15    : in     vl_logic;
        D0HSTXDATA14    : in     vl_logic;
        D0HSTXDATA13    : in     vl_logic;
        D0HSTXDATA12    : in     vl_logic;
        D0HSTXDATA11    : in     vl_logic;
        D0HSTXDATA10    : in     vl_logic;
        D0HSTXDATA9     : in     vl_logic;
        D0HSTXDATA8     : in     vl_logic;
        D0HSTXDATA7     : in     vl_logic;
        D0HSTXDATA6     : in     vl_logic;
        D0HSTXDATA5     : in     vl_logic;
        D0HSTXDATA4     : in     vl_logic;
        D0HSTXDATA3     : in     vl_logic;
        D0HSTXDATA2     : in     vl_logic;
        D0HSTXDATA1     : in     vl_logic;
        D0HSTXDATA0     : in     vl_logic;
        D0HSSEREN       : in     vl_logic;
        D0TXHSPD        : in     vl_logic;
        D0DRXHS         : out    vl_logic;
        D1DRXLPP        : out    vl_logic;
        D1RXLPEN        : in     vl_logic;
        D1DRXLPN        : out    vl_logic;
        D1DCDP          : out    vl_logic;
        D1CDEN          : in     vl_logic;
        D1DCDN          : out    vl_logic;
        D1DTXLPP        : in     vl_logic;
        D1TXLPEN        : in     vl_logic;
        D1DTXLPN        : in     vl_logic;
        D1RXHSEN        : in     vl_logic;
        D1HSRXDATA15    : out    vl_logic;
        D1HSRXDATA14    : out    vl_logic;
        D1HSRXDATA13    : out    vl_logic;
        D1HSRXDATA12    : out    vl_logic;
        D1HSRXDATA11    : out    vl_logic;
        D1HSRXDATA10    : out    vl_logic;
        D1HSRXDATA9     : out    vl_logic;
        D1HSRXDATA8     : out    vl_logic;
        D1HSRXDATA7     : out    vl_logic;
        D1HSRXDATA6     : out    vl_logic;
        D1HSRXDATA5     : out    vl_logic;
        D1HSRXDATA4     : out    vl_logic;
        D1HSRXDATA3     : out    vl_logic;
        D1HSRXDATA2     : out    vl_logic;
        D1HSRXDATA1     : out    vl_logic;
        D1HSRXDATA0     : out    vl_logic;
        D1SYNC          : out    vl_logic;
        D1ERRSYNC       : out    vl_logic;
        D1NOSYNC        : out    vl_logic;
        D1HSDESEREN     : in     vl_logic;
        D1TXHSEN        : in     vl_logic;
        D1HSTXDATA15    : in     vl_logic;
        D1HSTXDATA14    : in     vl_logic;
        D1HSTXDATA13    : in     vl_logic;
        D1HSTXDATA12    : in     vl_logic;
        D1HSTXDATA11    : in     vl_logic;
        D1HSTXDATA10    : in     vl_logic;
        D1HSTXDATA9     : in     vl_logic;
        D1HSTXDATA8     : in     vl_logic;
        D1HSTXDATA7     : in     vl_logic;
        D1HSTXDATA6     : in     vl_logic;
        D1HSTXDATA5     : in     vl_logic;
        D1HSTXDATA4     : in     vl_logic;
        D1HSTXDATA3     : in     vl_logic;
        D1HSTXDATA2     : in     vl_logic;
        D1HSTXDATA1     : in     vl_logic;
        D1HSTXDATA0     : in     vl_logic;
        D1HSSEREN       : in     vl_logic;
        D1TXHSPD        : in     vl_logic;
        D1DRXHS         : out    vl_logic;
        D2DRXLPP        : out    vl_logic;
        D2RXLPEN        : in     vl_logic;
        D2DRXLPN        : out    vl_logic;
        D2DCDP          : out    vl_logic;
        D2CDEN          : in     vl_logic;
        D2DCDN          : out    vl_logic;
        D2DTXLPP        : in     vl_logic;
        D2TXLPEN        : in     vl_logic;
        D2DTXLPN        : in     vl_logic;
        D2RXHSEN        : in     vl_logic;
        D2HSRXDATA15    : out    vl_logic;
        D2HSRXDATA14    : out    vl_logic;
        D2HSRXDATA13    : out    vl_logic;
        D2HSRXDATA12    : out    vl_logic;
        D2HSRXDATA11    : out    vl_logic;
        D2HSRXDATA10    : out    vl_logic;
        D2HSRXDATA9     : out    vl_logic;
        D2HSRXDATA8     : out    vl_logic;
        D2HSRXDATA7     : out    vl_logic;
        D2HSRXDATA6     : out    vl_logic;
        D2HSRXDATA5     : out    vl_logic;
        D2HSRXDATA4     : out    vl_logic;
        D2HSRXDATA3     : out    vl_logic;
        D2HSRXDATA2     : out    vl_logic;
        D2HSRXDATA1     : out    vl_logic;
        D2HSRXDATA0     : out    vl_logic;
        D2SYNC          : out    vl_logic;
        D2ERRSYNC       : out    vl_logic;
        D2NOSYNC        : out    vl_logic;
        D2HSDESEREN     : in     vl_logic;
        D2TXHSEN        : in     vl_logic;
        D2HSTXDATA15    : in     vl_logic;
        D2HSTXDATA14    : in     vl_logic;
        D2HSTXDATA13    : in     vl_logic;
        D2HSTXDATA12    : in     vl_logic;
        D2HSTXDATA11    : in     vl_logic;
        D2HSTXDATA10    : in     vl_logic;
        D2HSTXDATA9     : in     vl_logic;
        D2HSTXDATA8     : in     vl_logic;
        D2HSTXDATA7     : in     vl_logic;
        D2HSTXDATA6     : in     vl_logic;
        D2HSTXDATA5     : in     vl_logic;
        D2HSTXDATA4     : in     vl_logic;
        D2HSTXDATA3     : in     vl_logic;
        D2HSTXDATA2     : in     vl_logic;
        D2HSTXDATA1     : in     vl_logic;
        D2HSTXDATA0     : in     vl_logic;
        D2HSSEREN       : in     vl_logic;
        D2TXHSPD        : in     vl_logic;
        D2DRXHS         : out    vl_logic;
        D3DRXLPP        : out    vl_logic;
        D3RXLPEN        : in     vl_logic;
        D3DRXLPN        : out    vl_logic;
        D3DCDP          : out    vl_logic;
        D3CDEN          : in     vl_logic;
        D3DCDN          : out    vl_logic;
        D3DTXLPP        : in     vl_logic;
        D3TXLPEN        : in     vl_logic;
        D3DTXLPN        : in     vl_logic;
        D3RXHSEN        : in     vl_logic;
        D3HSRXDATA15    : out    vl_logic;
        D3HSRXDATA14    : out    vl_logic;
        D3HSRXDATA13    : out    vl_logic;
        D3HSRXDATA12    : out    vl_logic;
        D3HSRXDATA11    : out    vl_logic;
        D3HSRXDATA10    : out    vl_logic;
        D3HSRXDATA9     : out    vl_logic;
        D3HSRXDATA8     : out    vl_logic;
        D3HSRXDATA7     : out    vl_logic;
        D3HSRXDATA6     : out    vl_logic;
        D3HSRXDATA5     : out    vl_logic;
        D3HSRXDATA4     : out    vl_logic;
        D3HSRXDATA3     : out    vl_logic;
        D3HSRXDATA2     : out    vl_logic;
        D3HSRXDATA1     : out    vl_logic;
        D3HSRXDATA0     : out    vl_logic;
        D3SYNC          : out    vl_logic;
        D3ERRSYNC       : out    vl_logic;
        D3NOSYNC        : out    vl_logic;
        D3HSDESEREN     : in     vl_logic;
        D3TXHSEN        : in     vl_logic;
        D3HSTXDATA15    : in     vl_logic;
        D3HSTXDATA14    : in     vl_logic;
        D3HSTXDATA13    : in     vl_logic;
        D3HSTXDATA12    : in     vl_logic;
        D3HSTXDATA11    : in     vl_logic;
        D3HSTXDATA10    : in     vl_logic;
        D3HSTXDATA9     : in     vl_logic;
        D3HSTXDATA8     : in     vl_logic;
        D3HSTXDATA7     : in     vl_logic;
        D3HSTXDATA6     : in     vl_logic;
        D3HSTXDATA5     : in     vl_logic;
        D3HSTXDATA4     : in     vl_logic;
        D3HSTXDATA3     : in     vl_logic;
        D3HSTXDATA2     : in     vl_logic;
        D3HSTXDATA1     : in     vl_logic;
        D3HSTXDATA0     : in     vl_logic;
        D3HSSEREN       : in     vl_logic;
        D3TXHSPD        : in     vl_logic;
        D3DRXHS         : out    vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of HSEL : constant is 1;
    attribute mti_svvh_generic_type of HS_16BIT_EN : constant is 1;
    attribute mti_svvh_generic_type of CN : constant is 1;
    attribute mti_svvh_generic_type of CM : constant is 1;
    attribute mti_svvh_generic_type of CO : constant is 1;
    attribute mti_svvh_generic_type of PLL_TST : constant is 1;
    attribute mti_svvh_generic_type of ENP_DESER : constant is 1;
end MIPIDPHYA;
