library verilog;
use verilog.vl_types.all;
entity config_sspi_inst_dec is
    port(
        sspi_async_rst  : in     vl_logic;
        clk             : in     vl_logic;
        instruction     : in     vl_logic_vector(7 downto 0);
        sspi_xflash     : in     vl_logic;
        sspi_xsram      : in     vl_logic;
        sspi_idle       : in     vl_logic;
        cmd_inf_r       : in     vl_logic;
        csspi           : in     vl_logic;
        decrypt_en      : in     vl_logic;
        prgincr_int_ctrl: in     vl_logic;
        addrshift_o     : out    vl_logic;
        inc_inst        : out    vl_logic;
        progdis_o       : out    vl_logic;
        rst_addr_o      : out    vl_logic;
        xprogen_ee_o    : out    vl_logic;
        xreaden_sram_o  : out    vl_logic;
        erase_tag_o     : out    vl_logic;
        erase_ee_o      : out    vl_logic;
        eraseall_ee_o   : out    vl_logic;
        sspi_erase      : out    vl_logic;
        sspi_read_en_ee : out    vl_logic;
        sram_read       : out    vl_logic;
        flash_read      : out    vl_logic;
        vfy_reg32_inst  : out    vl_logic;
        read_o          : out    vl_logic;
        vfy_incr_o      : out    vl_logic;
        ucode_o         : out    vl_logic;
        ucode_ee_o      : out    vl_logic;
        idcode_o        : out    vl_logic;
        read_ee_o       : out    vl_logic;
        read_tag_o      : out    vl_logic;
        prog_tag_o      : out    vl_logic;
        progstatus_ee_o : out    vl_logic;
        readstatus_ee_o : out    vl_logic;
        prog_inc_ee_o   : out    vl_logic;
        progenc_inc_ee_o: out    vl_logic;
        progucode_ee_o  : out    vl_logic;
        progsec_ee_o    : out    vl_logic;
        progdone_ee_o   : out    vl_logic;
        vfy_incr_ee_o   : out    vl_logic;
        progctrl0_ee_o  : out    vl_logic;
        vfyctrl0_ee_o   : out    vl_logic;
        vfyctrl0_o      : out    vl_logic;
        refresh_o       : out    vl_logic;
        progcrc32_ee_o  : out    vl_logic;
        vfycrc32_o      : out    vl_logic;
        vfycrc32_ee_o   : out    vl_logic;
        selasr          : out    vl_logic;
        seldsr          : out    vl_logic;
        sspi_fl_ep      : out    vl_logic;
        sspi_fl_ep_only : out    vl_logic;
        prog_inst       : out    vl_logic;
        vfy_inst        : out    vl_logic;
        protect_shift_o : out    vl_logic;
        rst_flash_status: out    vl_logic;
        rst_16_crc_r    : out    vl_logic;
        read_16_crc     : out    vl_logic;
        progenc_inc_flash: out    vl_logic;
        sspi_refresh_r  : out    vl_logic
    );
end config_sspi_inst_dec;
