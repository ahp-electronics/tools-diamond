--
@ER--RbBF$osHE50RO42RgRgg1b$MDHHO0R$,Q3MO
R--RDqDRosHER0#sCC#s8PC3-
-
R--fN]C8:CsR#//$DMbH0OH$N/lb..jjDjdNl0/NCbbsO#/b/D8D/HLo_CMD0N0H/OCN388PyE84
Rf-
-
---
-CRoMNCs0bCRsNFboCN0RDOCDO3RNkDODCN0#NROsCsH#NRL#RC8FoMRCbM/sRFbHkMb0-#
-H
DLssN$CRHC
C;kR#CHCCC38#0_oDFH4O_43ncN;DD
0CMHR0$oDb_CRNVH
#RSMoCCOsHRS5
Sx#HCRR:HCM0oRCs:4=R
;S2
FSbs50R
oSSCkMF0RR:FRk0#_08DHFoOS;
SFbsb0FkRF:Rk#0R0D8_FOoH;S
SO0FkRF:Rk#0R0D8_FOoH_OPC05Fs#CHx-84RF0IMF2Rj;S
SoHCMMRR:H#MR0D8_FOoH_OPC05Fs#CHx-84RF0IMF2Rj;S
SbbsFH:MRRRHM#_08DHFoOC_POs0F5x#HCR-48MFI0jFR2S;
SMOHRH:RM0R#8F_Do2HO;M
C8bRo_NDCV
;
NEsOHO0C0CksRFLFDMCNRRFVoDb_CRNVH
#RSo#HMRND0Ro:#_08DHFoOC_POs0F5x#HCR-48MFI0jFR2S;
#MHoN0DRb#:R0D8_FOoH_OPC05Fs#CHx-84RF0IMF2Rj;C
Lo
HMS50bj<2R=sRbFMbH5;j2
oS05Rj2<o=RCMMH5;j2
FSOkj052=R<R50ojF2Rs0R5b25jR8NMRMOH2
;SSFbsO#C#RH5OMb,RsHFbMo,RCMMH,oR0,bR02SR
SsPNHDNLCRRH:MRH0CCosS;
LHCoMS
SVRFsHMRHR04RFHR#x4C-RFDFbS
SS50bH<2R=sRbFMbH5RH2NRM80Hb5-;42
SSS0Ho52=R<RMoCHHM52sRFRs5bFMbH5RH2NRM80Ho5-242;S
SSkOF025HRR<=0Ho52sRFRb505RH2NRM8O2HM;S
SCRM8DbFF;C
SMb8RsCFO#
#;SMoCFRk0<0=RoH5#x4C-2S;
bbsFFRk0<0=RbH5#x4C-2
;
CRM8LDFFC;NM
-
-
R--OsNs$FRDFE	NCRN8NC88sHRI00ERIDFRCDPC#VRFRFDF	ERNC
N8-H-RMs0ClHC8NR0CNC88sN#RssCRHDbbC8RN8#Cs

--DsHLNRs$HCCC;#
kCCRHC#C30D8_FOoH_n44cD3NDC;
M00H$8RN8bsoR
H#SMoCCOsHRS5
Sx#HCRR:HCM0oRCs:.=RgS;
SNDCVx#HCRR:HCM0oRCs:n=R
;S2
FSbs50R
OSSFRk0:kRF00R#8F_Do;HO
8SSRF:Rk#0R0D8_FOoH_OPC05Fs#CHx-84RF0IMF2Rj;S
SNRR:H#MR0D8_FOoH_OPC05Fs#CHx-84RF0IMF2Rj;S
SLRR:H#MR0D8_FOoH_OPC05Fs#CHx-84RF0IMF2Rj;S
SORHM:MRHR8#0_oDFH;O2
8CMR8N8s;ob
s
NO0EHCkO0sLCRFCFDNFMRV8RN8bsoR
H#
kSVMHO0FOMRNODOM50RO#FM00NMR,#xRNDCVR#x:MRH0CCoss2RCs0kMMRH0CCos#RH
NSPsLHNDDCRC0NVlsb,ORM0:MRH0CCosS;
LHCoMS
SDVCN0Rlb:#=RxRR/DVCN#
x;SVSHR#55xFRl8CRDNxV#2RR=j02RE
CMSsSSORM0:D=RC0NVl;bR
CSSDR#C
SSSs0OMRR:=5NDCVb0lR4+R2S;
S8CMR;HV
sSSCs0kMORsM
0;S8CMRDONO0OM;S

O#FM00NMRNDCV0OMRH:RMo0CC:sR=NRODMOO0H5#xRC,DVCN#CHx2
;
SMVkOF0HMER0HC#DNHV#x5CRO#FM00NMR:MRR0HMCsoC2CRs0MksR0HMCsoCR
H#SsPNHDNLCxR#RH:RMo0CC
s;SoLCHSM
SRHV5=MRRC5DNMVO02-42ER0C
MRS#SSx=R:Rx#HCFRl8CRDNHV#x
C;SHSSV#R5xRR=j02RERCM
SSSSR#x:D=RC#NVH;xCRS
SS8CMR;HV
CSSD
#CS#SSx=R:RNDCVx#HCS;
S8CMR;HV
sSSCs0kMxR#;C
SM08REDH#C#NVH;xC
V
Sk0MOHRFMlLNGH50RO#FM00NMR:MRR0HMCsoC2CRs0MksR0HMCsoCR
H#SsPNHDNLCNRlGRR:HCM0o;Cs
CSLo
HMSNSlG=R:R+5M4D2*C#NVHRxC-;R4
HSSVlR5N>GR=HR#xRC20MEC
SSSlRNG:#=RH-xC4S;
S8CMR;HV
sSSCs0kMNRlGS;
CRM8lLNGH
0;
HS#oDMNRMoCNRL:#_08DHFoOC_POs0F5x#HCR-48MFI0jFR2S;
#MHoNbDRsNFbL#:R0D8_FOoH_OPC05Fs#CHx-84RF0IMF2Rj;#
SHNoMDHROMR0:#_08DHFoOC_POs0F5NDCV0OMRI8FMR0Fj
2;So#HMRNDO0HML#:R0D8_FOoH_OPC05FsDVCNORM08MFI0jFR2S;
#MHoNODRs0HM:0R#8F_Do_HOP0COF#s5HRxC8MFI0jFR2S;
#MHoNoDRCkMF0RR:#_08DHFoOS;
#MHoNbDRsFFbk:0RR8#0_oDFH
O;
FSOlMbFCRM0oDb_CRNVH
#RSCSoMHCsO
R5S#SSHRxC:MRH0CCosS
S2S;
SsbF0
R5SoSSCkMF0RR:FRk0#_08DHFoOS;
SsSbFkbF0RR:FRk0#_08DHFoOS;
SFSOk:0RR0FkR8#0_oDFHPO_CFO0sH5#x4C-RI8FMR0Fj
2;SoSSCMMHRH:RM0R#8F_Do_HOP0COF#s5H-xC4FR8IFM0R;j2
SSSbbsFH:MRRRHM#_08DHFoOC_POs0F5x#HCR-48MFI0jFR2S;
SHSOMRR:H#MR0D8_FOoH2S;
CRM8ObFlFMMC0
;
SlOFbCFMMN0R8H8sbCbDR
H#SCSoMHCsO
R5S#SSHRxC:MRH0CCosS
S2S;
SsbF0
R5SOSSFRk0:kRF00R#8F_Do;HO
SSS8RR:FRk0#_08DHFoOC_POs0F5x#HCR-48MFI0jFR2S;
SRSN:MRHR8#0_oDFHPO_CFO0sH5#x4C-RI8FMR0Fj
2;SLSSRH:RM0R#8F_Do_HOP0COF#s5H-xC4FR8IFM0R;j2
SSSORHM:MRHR8#0_oDFHSO
S
2;S8CMRlOFbCFMM
0;
FSOlMbFCRM0BAYuzHwR#SR
SsbF0
R5SRSN:MRHR8#0_oDFH
O;SRSL:kRF00R#8F_Do
HOS;S2
MSC8FROlMbFC;M0
#
SHNoMDoRL,RLb:0R#8F_Do_HOP0COF#s5H-xC4FR8IFM0R;j2
HS#oDMNR0Lo,0LbR#:R0D8_FOoH_OPC05Fs#CHx-84RF0IMF2Rj;#
SHNoMD,RobRR:#_08DHFoOC_POs0F5NDCV0OM-84RF0IMF2Rj;#
SHNoMDLRo,RbL:0R#8F_Do_HOP0COFDs5CONVM40-RI8FMR0Fj
2;So#HMRNDVRFF:0R#8F_Do;HO
oLCH
M
SMoCN<LR=RRNNRM8LS;
bbsFN<LR=RRNFLsR;O
SH5M0j<2R=HROMS;
O0HML25jRR<=O;HM
-
S-CR	C0bREDCRNDLC#ER#FRs0F0sREMCRN#lCR0oCRF0FRMDFoq
S:FRVsRRMHjMRRR0FDVCNO-M04CRoMNCs0SC
SMOF#M0N0GRlL:0RR0HMCsoCRR:=lLNGHM052S;
SMOF#M0N0VRD#:xRR0HMCsoCRR:=0#EHDVCN#CHx5;M2
OSSF0M#NRM0l0MLRH:RMo0CC:sR=CRDNHV#xMC*;S
SO#FM00NMRDNDF#MCR#:R0D8_FOoH_OPC05Fsl0GLRI8FMR0Fl0ML2=R:R05FE#Cs='>R4;'2
CSLoRHM
LSSoM5lLR02<o=RCLMN5LlM0
2;SbSL5LlM0<2R=sRbFLbN5LlM0
2;SoSL0M5lLR02<L=RoM5lL;02
LSSbl05M2L0RR<=Llb5M2L0;S

SR--OONDk0DNCER0CHRL0H-I#oCR'N#RMb8R'N#RML8RkCVVsER0CSl
SRA:VRFslMRHRLlM0R+40lFRGRL0oCCMsCN0RS
SS0Lo5Rl2<o=RCLMN5Rl2F5sRbbsFNlL52MRN8oRL0-5l4;22
SSSA:tXRuBYARzwb0FsRblNRo5L025l,oRL52l2;S
SS0Lb5Rl2<b=RsNFbL25lR8NMR0Lb54l-2S;
SuSAXB:RYzuAwFRbsl0RN5bRL5b0lR2,Llb52
2;SMSC8CRoMNCs0
C;
-SS-FROb0$REDCRC'NV#RRoNRM8bsRVF0lRELCRoMRN8bRL
oSSL25MRR<=Llo5G2L0;S
SbML52=R<R5Lbl0GL2
;
S-S-RVLkVRCs0RECOsNs$MRHRs5VF0lREOCRN$ssRMoCC0sNFRs2
BSS:VRHRR5M/j=R2CRoMNCs0
CRSBSSARX:BAYuzbwRFRs0l5NbO0HM5,M2RMOH0ML52
2;SMSC8CRoMNCs0
C;
-SS-NRODDOkNR0C0RECL-H0ICH#RsONs#HCRFVslER0CHRL0H-I#oCRbR'#NRM8O
HMS:S8RRHV5LlG0RR>l0ML2CRoMNCs0
CRSCSS:FRVsRRlHlMRGRL08MFI0lFRM+L04CRoMNCs0SC
SOSSs0HM5Rl2<L=Ro-5l4F2RsOR5HLM05RM2NRM8Llb5-242;S
SS8CMRMoCC0sNCS;
S8CMRMoCC0sNCS;
SHOsMl05M2L0RR<=O0HML25M;S

SR--OONDk0DNCER0CkR#lS
S8G5lL80RF0IMFMRlLR02<N=R5LlG0FR8IFM0RLlM0S2
SFSGs5RLl0GLRI8FMR0Fl0ML2FRGssROH5M0l0GLRI8FMR0Fl0ML2S;
CRM8oCCMsCN0;S

-o-RCsMCNR0C0RECOsNsH
C#S:OoR_obDVCN
oSSCsMCHlORN5bR
SSS#CHxRR=>DVCNO
M0S
S2SFSbsl0RN5bR
SSSoFCMk=0R>CRoM0Fk,S
SSFbsb0FkRR=>bbsFF,k0
SSSO0FkRR=>O0HM5NDCV0OMRI8FMR0F4
2,SoSSCMMHRR=>oDL5CONVM40-RI8FMR0Fj
2,SbSSsHFbM>R=R5bLDVCNO-M04FR8IFM0R,j2
SSSORHM=O>RHSM
S
2;
FSOk<0R=HROMD05CONVM;02
M
C8FRLFNDCM
;
---
-kRVDsDRHDbbC8RN8
Cs-D-
HNLssH$RC;CC
Ck#RCHCC03#8F_Do_HO4c4n3DND;M
C0$H0R8N8sbHbDHCR#o
SCsMCH5OR
#SSHRxC:MRH0CCos=R:RSg
2S;
b0FsRS5
SkOF0RR:FRk0#_08DHFoOS;
S:8RR0FkR8#0_oDFHPO_CFO0sH5#x4C-RI8FMR0Fj
2;SRSN:MRHR8#0_oDFHPO_CFO0sH5#x4C-RI8FMR0Fj
2;SRSL:MRHR8#0_oDFHPO_CFO0sH5#x4C-RI8FMR0Fj
2;SHSOMRR:H#MR0D8_FOoH2C;
MN8R8H8sbCbD;N

sHOE00COkRsCLDFFCRNMFNVR8H8sbCbDR
H#So#HMRNDoFCMk:0RR8#0_oDFH
O;So#HMRNDbbsFFRk0:0R#8F_Do;HO
HS#oDMNRMOH0#:R0D8_FOoH_OPC05Fs#CHxRI8FMR0Fj
2;So#HMRNDoNCML#:R0D8_FOoH_OPC05Fs#CHx-84RF0IMF2Rj;#
SHNoMDsRbFLbN:0R#8F_Do_HOP0COF#s5H-xC4FR8IFM0R;j2
oLCHSM
oNCML=R<RNNRML8R;b
SsNFbL=R<RFNRs;RL
HSOM#05HRxC8MFI04FR2=R<Rs5bFLbNR8NMRMOH0H5#x4C-RI8FMR0FjR22FosRCLMN;O
SH5M0j<2R=HROMS;
8=R<RGNRFLsRRsGFRMOH0H5#x4C-RI8FMR0Fj
2;SkOF0=R<RMOH0H5#x;C2
8CMRFLFDMCN;-

--
-Rb0FRPDCCCDRM00H$FRVs8RN8RCsoCCMsFN0s-
-RCk##HRsbCbDRRHVD#C#RN0EMqRvXu)Qu,p R#CDC#RkCO#RN$ssRFDF	CNEN-8
-H
DLssN$CRHCRC;
Ck#RCHCC03#8F_Do_HO4c4n3DND;M
C0$H0R7q7R
H#RRRRoCCMs5HOI0H8ERR:HCM0oRCs:4=RnR2;-[-RNRo
RbRRF5s0qH:RM0R#8F_Do_HOP0COFIs5HE80RR-48MFI0jFR2R;
RRRRRRRRAH:RM0R#8F_Do_HOP0COFIs5HE80RR-48MFI0jFR2R;
RRRRRRRRBRQh:MRHR8#0_oDFH
O;RRRRRRRRR:mRR0FkR8#0_oDFHPO_CFO0sH5I8R0E-84RF0IMF2Rj;R
RRRRRRBRRm:zaR0FkR8#0_oDFH;O2
8CMR7q7;N

sHOE00COkRsCODCD_PDCCFDRV7Rq7#RH
FSOMN#0Mv0RqQX)u upRH:RMo0CC:sR=;RU
V
Sk0MOHRFMOONDDVCN#CHxRF5OMN#0MI0R:MRH0CCoss2RCs0kMMRH0CCos#RH
PSSNNsHLRDCsDPN:0HMCsoCRR:=4S;
LHCoMS
SIDEHCsR5PRND*PRsN<DRRRI2DbFF
SSSsDPNRR:=sDPNR4+R;S
SCRM8DbFF;S
SH5VRsDPNRc<R2ER0C
MRSsSSPRND:c=R;SR
S8CMR;HV
sSSCs0kMPRsN
D;S8CMRDONONDCVx#HC
;
SlOFbCFMMN0R8o8sb#RH
oSSCsMCH5OR
SSS#CHxRH:RMo0CC
s;SDSSC#NVHRxC:MRH0CCosSR
S
2;SFSbs50R
SSSO0FkRF:Rk#0R0D8_FOoH;S
SS:8RR0FkR8#0_oDFHPO_CFO0sH5#x4C-RI8FMR0Fj
2;SNSSRH:RM0R#8F_Do_HOP0COF#s5H-xC4FR8IFM0R;j2
SSSLRR:H#MR0D8_FOoH_OPC05Fs#CHx-84RF0IMF2Rj;S
SSMOHRH:RM0R#8F_Do
HOS;S2
MSC8FROlMbFC;M0
O
SFFlbM0CMR8N8sbHbDHCR#S
SoCCMsRHO5S
SSx#HCRR:HCM0o
CsS;S2
bSSFRs05S
SSkOF0RR:FRk0#_08DHFoOS;
SRS8:kRF00R#8F_Do_HOP0COF#s5H-xC4FR8IFM0R;j2
SSSNRR:H#MR0D8_FOoH_OPC05Fs#CHx-84RF0IMF2Rj;S
SS:LRRRHM#_08DHFoOC_POs0F5x#HCR-48MFI0jFR2S;
SHSOMRR:H#MR0D8_FOoH
2SS;C
SMO8RFFlbM0CM;L

CMoH
NSL:VRHRH5I8R0E>qRvXu)Qu2p RMoCC0sNCS
SNR4:Ns88o
bRSoSSCsMCHlORN5bR
SSSSx#HC>R=R8IH0
E,SSSS-D-RC#NVHRxC=O>RNDDOC#NVH5xCI0H8ES2
SDSSC#NVHRxC=c>R
SSS2S
SSsbF0NRlb
R5SSSSO0FkRR=>O0Fk,S
SSRS8=F>R,S
SSRSN=N>R,S
SSRSL=L>R,S
SSHSOM>R=RMOH
SSS2S;
CRM8oCCMsCN0;S

#RN:H5VRI0H8E=R<RXvq)uQupR 2oCCMsCN0
NSS4N:R8H8sbCbDRS
SSMoCCOsHRblNRS5
S#SSHRxC=I>RHE80
SSS2S
SSsbF0NRlb
R5SSSSO0FkRR=>O0Fk,S
SSRS8=F>R,S
SSRSN=N>R,S
SSRSL=L>R,S
SSHSOM>R=RMOH
SSS2S;
CRM8oCCMsCN0;C

MO8RC_DDDCCPD
;

