library verilog;
use verilog.vl_types.all;
entity MPC_TOP is
    port(
        MC1_PAR_ODD     : in     vl_logic;
        MPI_PAR_CHK     : in     vl_logic;
        MPI_DP_ENABLE   : in     vl_logic;
        MPI_DMA_ENABLE  : in     vl_logic;
        DMA_TA          : in     vl_logic;
        DMA_RETRY       : in     vl_logic;
        DMA_TEA         : in     vl_logic;
        DMA_TRI_DATA    : in     vl_logic;
        DMA_TRI_CTL     : in     vl_logic;
        DMA_RD_DATA     : in     vl_logic_vector(0 to 31);
        DMA_RD_PARITY   : in     vl_logic_vector(0 to 3);
        MPC_CLK         : in     vl_logic;
        MPC_TSIZ        : in     vl_logic_vector(0 to 1);
        MPC_READ        : in     vl_logic;
        MPC_BURST       : in     vl_logic;
        MPC_BDIP        : in     vl_logic;
        MPC_TS          : in     vl_logic;
        MPC_ADDR        : in     vl_logic_vector(14 to 31);
        MPC_CS0         : in     vl_logic;
        MPC_CS1         : in     vl_logic;
        MPC_TA          : out    vl_logic;
        MPC_RETRY       : out    vl_logic;
        MPC_TEA         : out    vl_logic;
        MPC_TRI_DATA    : out    vl_logic;
        MPC_TRI_CTL     : out    vl_logic;
        MPC_WR_DATA     : in     vl_logic_vector(0 to 31);
        MPC_RD_DATA     : out    vl_logic_vector(0 to 31);
        MPC_WR_PARITY   : in     vl_logic_vector(0 to 3);
        MPC_RD_PARITY   : out    vl_logic_vector(0 to 3);
        MPC_RESET_N     : in     vl_logic;
        AHB_RESET_N     : in     vl_logic;
        BUS_SIZE        : in     vl_logic_vector(2 downto 0);
        MPC_SYNC        : in     vl_logic;
        HCLK            : in     vl_logic;
        AHB_BUS_GNT     : in     vl_logic;
        AHB_READY       : in     vl_logic;
        AHB_RD_DATA     : in     vl_logic_vector(31 downto 0);
        AHB_RD_PARITY   : in     vl_logic_vector(3 downto 0);
        AHB_RESP        : in     vl_logic_vector(1 downto 0);
        AHB_BUS_REQ     : out    vl_logic;
        AHB_BUS_LOCK    : out    vl_logic;
        AHB_BURST       : out    vl_logic;
        AHB_SIZE        : out    vl_logic_vector(1 downto 0);
        AHB_WRITE       : out    vl_logic;
        AHB_ADDR        : out    vl_logic_vector(17 downto 0);
        AHB_IRQ         : out    vl_logic;
        AHB_TRANS       : out    vl_logic_vector(1 downto 0);
        AHB_WR_DATA     : out    vl_logic_vector(31 downto 0);
        AHB_WR_PARITY   : out    vl_logic_vector(3 downto 0);
        SCANEN          : in     vl_logic
    );
end MPC_TOP;
