library verilog;
use verilog.vl_types.all;
entity ctl_spare_gate is
    port(
        signal_in       : in     vl_logic
    );
end ctl_spare_gate;
