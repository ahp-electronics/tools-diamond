library verilog;
use verilog.vl_types.all;
entity vlom4mce is
    port(
        Z               : out    vl_logic
    );
end vlom4mce;
