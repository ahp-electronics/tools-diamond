library verilog;
use verilog.vl_types.all;
entity cfg_front is
    generic(
        MASTER_SERI     : integer := 8;
        MASTER_PARA     : integer := 12;
        ASYNC_PERI      : integer := 13;
        SLAVE_SERI      : integer := 15;
        SLAVE_PARA      : integer := 9;
        FPSC_PARA       : integer := 7;
        MASTER_BYTE     : integer := 6;
        FLASH_SPI03     : integer := 5;
        FLASH_SPIX      : integer := 4;
        MPC_BYTE        : integer := 10;
        MPC_HWORD       : integer := 11;
        MPC_WORD        : integer := 14;
        CHK_PRE         : integer := 0;
        CHK_ID          : integer := 1;
        CHK_HDR         : integer := 2;
        CHK_FPGA        : integer := 3;
        CHK_RAM         : integer := 6;
        CHK_FPSC        : integer := 5;
        CHK_POST        : integer := 7
    );
    port(
        CODE0           : in     vl_logic_vector(7 downto 0);
        CODE1           : in     vl_logic_vector(7 downto 0);
        CODE2           : in     vl_logic_vector(7 downto 0);
        CODE3           : in     vl_logic_vector(7 downto 0);
        CODE4           : in     vl_logic_vector(7 downto 0);
        CODE5           : in     vl_logic_vector(7 downto 0);
        CODE6           : in     vl_logic_vector(7 downto 0);
        CODE7           : in     vl_logic_vector(7 downto 0);
        IDCODE3         : in     vl_logic_vector(7 downto 0);
        IDCODE4         : in     vl_logic_vector(7 downto 0);
        IDCODE5         : in     vl_logic_vector(7 downto 0);
        IDCODE6         : in     vl_logic_vector(7 downto 0);
        IDCODE7         : in     vl_logic_vector(7 downto 0);
        J_SPI_PROG      : in     vl_logic;
        J_SHDR          : in     vl_logic;
        J_SCANIN        : in     vl_logic;
        J_TCK           : in     vl_logic;
        RCLKS           : in     vl_logic;
        CCLK            : in     vl_logic;
        SER_CCLK        : in     vl_logic;
        CFRONT_INIT_N   : in     vl_logic;
        DEC_EN          : in     vl_logic;
        CS0_N           : in     vl_logic;
        CS1             : in     vl_logic;
        WR_N            : in     vl_logic;
        MODE            : in     vl_logic_vector(3 downto 0);
        PRGM_JTAG       : in     vl_logic;
        PRGM_SYS        : in     vl_logic_vector(2 downto 0);
        MPI_CLK_RAM     : in     vl_logic;
        FPSC_CLK_RAM    : in     vl_logic;
        USR_CLK_RAM     : in     vl_logic;
        OSC_CLK_RAM     : in     vl_logic;
        DIS_MODES_RAM   : in     vl_logic;
        EXT_CCLK_RAM    : in     vl_logic;
        TEST_CTR_RAM    : in     vl_logic;
        RST_BUS_RAM_N   : in     vl_logic;
        RST_HCLK_RAM_N  : in     vl_logic;
        RST_RAM_RAM_N   : in     vl_logic;
        EN_MPI_PARITY_RAM: in     vl_logic;
        MODE_RAM        : in     vl_logic_vector(3 downto 0);
        STRT_RAM        : in     vl_logic_vector(4 downto 0);
        TRI_RAM         : in     vl_logic_vector(3 downto 0);
        SPI_ADDR_RAM    : in     vl_logic_vector(31 downto 0);
        SYS_DATA_RDY    : in     vl_logic;
        SYS_CFGD_BYTE   : in     vl_logic_vector(7 downto 0);
        DEL_D           : in     vl_logic_vector(7 downto 0);
        DONE            : in     vl_logic;
        PAD_INIT_N      : in     vl_logic;
        PWR_ON          : in     vl_logic;
        SERIAL_DATA     : in     vl_logic;
        SYS_DAISY       : in     vl_logic;
        MPI_USR_ENABLE  : in     vl_logic;
        RD_CFG_JTAG     : in     vl_logic;
        TDI_JTAG        : in     vl_logic;
        BS_MODE         : in     vl_logic;
        SYS_MODE        : in     vl_logic;
        CHK_STATE       : in     vl_logic_vector(2 downto 0);
        READ_START      : in     vl_logic;
        HDC             : out    vl_logic;
        LDC_N           : out    vl_logic;
        CFGDOUT_JTAG_N  : out    vl_logic;
        M_CFRONT_INIT_N : out    vl_logic;
        RDY_BUSY_N      : out    vl_logic;
        DOUT            : out    vl_logic;
        QOUT            : out    vl_logic;
        PRDY_TS         : out    vl_logic;
        PA_OUT          : out    vl_logic_vector(21 downto 0);
        ADDR_TS         : out    vl_logic;
        EN_CCLK_N       : out    vl_logic;
        MPI_DP_ENABLE   : out    vl_logic;
        RST_BUS         : out    vl_logic;
        HCLK_RST        : out    vl_logic;
        CLKMPI          : out    vl_logic;
        CLKFPSC         : out    vl_logic;
        CLKUSR          : out    vl_logic;
        CLKOSC          : out    vl_logic;
        EXTCCLK         : out    vl_logic;
        GSRNRAM         : out    vl_logic;
        TRIRAM          : out    vl_logic;
        RSTRAM          : out    vl_logic;
        DEL_D_REG       : out    vl_logic_vector(7 downto 0);
        P2S_REG0        : out    vl_logic;
        SYS_BUS_DEC     : out    vl_logic;
        MASTER_SERI_DEC_REG: out    vl_logic;
        SYS_P2S_DONE    : out    vl_logic;
        STOPCCLK_N      : out    vl_logic;
        SYS_BUS_CFG     : out    vl_logic;
        LMODE           : out    vl_logic_vector(3 downto 0);
        M_CLK           : out    vl_logic
    );
end cfg_front;
