--
@ER--B$FbsEHo0OR52gR4g-cRRj.jd$R1MHbDO$H0ROQM
R--fN]C8:CsR#//$DMbH0OH$N/lb..jjDjdNl0/NCbbsN#/0D0/HoL/CFM_scONCN/sl__sIE3P8Ry4f-
-
-

--
-
R--7DkN-sbF0qR)vHRI0#ERCsbCNR0Cq)77 R11VRFss8CNR8NMRHIs0-C
-NRas0oCRp:RkMOC0RR-mq)BR
dB-D-
HNLssH$RC;CC
Ck#RCHCC03#8F_Do_HO4c4n3DND;#
kCCRHC#C30D8_FOoH_o#HM3C8N;DD
Ck#RCHCC03#8F_Do_HON0sHED3NDD;
HNLssF$RsdON;#
kCsRFO3NdFNsOObFl3DND;M
C0$H0Rv)q_W)_R
H#RRRRoCCMsRHO5R
RRRRRRNRVl$HD:0R#soHMRR:="MMFC
";RRRRRRRRI0H8ERR:HCM0oRCs:(=R;RR
RRRRRNRR8I8sHE80RH:RMo0CC:sR=;R(RRRRRRRR-L-RHCoRMoFkEFRVsCR8b
0ERRRRRRRR80CbERR:HCM0oRCs:R=R4;.U
RRRRRRRRk8F0C_soRR:LDFFCRNM:V=RNCD#;RRRR-R-R#ENR0FkbRk0s
CoRRRRRRRR8_HMsRCo:FRLFNDCM=R:RDVN#RC;RRRRRR--ERN#8NN0RbHMks0RCRo
RRRRRsRRNs88_osCRL:RFCFDN:MR=NRVD;#CRRRR-E-RNs8RCRN8Ns88CR##s
CoRRRRRRRRI8N8sC_soRR:LDFFCRNM:V=RNCD#RRRRRR--ERN8I0sHC8RN8#sC#CRsoR
RRRRRR;R2
RRRRsbF0
R5RRRRRRRR7amzRRR:FRk0#_08DHFoOC_POs0F58IH04E-RI8FMR0Fj
2;RRRRRRRR)7q7)RR:HRMR#_08DHFoOC_POs0F58N8s8IH04E-RI8FMR0Fj
2;RRRRRRRR7RQhRRR:HRMR#_08DHFoOC_POs0F58IH04E-RI8FMR0Fj
2;RRRRRRRRW7q7)RR:HRMR#_08DHFoOC_POs0F58N8s8IH04E-RI8FMR0Fj
2;RRRRRRRRWR RRRR:HRMR#_08DHFoOR;RRRRRRR--I0sHCMRCNCLDRsVFRlsN
RRRRRRRRiBpR:RRRRHMR8#0_oDFHRO;RRRRR-R-RFODOV	RFssRNRl,Ns88,HR8MR
RRRRRRBRmpRiR:MRHR0R#8F_DoRHORRRRR-RR-bRF0DROFRO	VRFs80Fk
RRRRRRRR
2;CRM8CHM00)$Rq)v__
W;

---w-RH0s#RbHlDCClM00NHRFMl0k#RRLCODNDCN8RsjOE

--NEsOHO0C0CksRONsEFjRVqR)v__)W#RH
MOF#M0N0kRMlC_OD_D#8bCCRH:RMo0CC:sR=5R580CbERR-4d2/.R2;RRRRRRRR-y-RRRFVs#FIRRFV7dB .RXcODCD#CRMC88C
MOF#M0N0kRMlC_OD_D#ICH8RH:RMo0CC:sR=5R5I0H8ERR-4c2/2R;RRRRRRRRR-y-RRRFVOkFDlRM#F7VRB. dXOcRC#DDRCMC8
C80C$bR0Fk_#Lk_b0$C#RHRsNsN5$RM_klODCD#C_8C8bRF0IMF,RjRk5MlC_OD_D#ICH8*+c2dFR8IFM0RRj2F#VR0D8_FOoH;H
#oDMNR0Fk_#LkRF:RkL0_k0#_$;bCRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--.N7Rs$sNRRFV80FkRM5HbRk000FRs#H-0CN0##2
HNoMDkRF0M_CRRRR:0R#8F_Do_HOP0COFMs5kOl_C#DD_C8CbFR8IFM0R;j2R-R-RNCML#DCRsVFRH0s-N#00
C##MHoNIDRb_CjCRMRR#:R0D8_FOoH_OPC05FsM_klODCD#C_8C8bRF0IMF2Rj;-RR-sRIHR0CCLMNDRC#VRFsCENORIsFRRFV)RqvODCD#H
#oDMNRCIb4M_CR:RRR8#0_oDFHPO_CFO0sk5MlC_OD_D#8bCCRI8FMR0FjR2;RR--I0sHCMRCNCLD#FRVsNRCOsERFFIRVqR)vCROD
D##MHoNHDRMC_soRRRR#:R0D8_FOoH_OPC05FsI0H8ER+d8MFI0jFR2R;RRRRRR-RR-#RkC08RFCRso0H#C7sRQ
hR#MHoNWDR  _)tR4RR#:R0D8_FOoH;H
#oDMNR_HMs4CoR:RRR8#0_oDFHPO_CFO0sH5I8+0EdFR8IFM0R;j2RRRR
o#HMRNDF_k0sRCoRRR:#_08DHFoOC_POs0F58IH0dE+RI8FMR0FjR2;RRRRRRRR-k-R#RC80sFRC#oH0RCs7amz
o#HMRNDs_N8sRCoRRR:#_08DHFoOC_POs0F58N8s8IH04E-RI8FMR0FjR2;RRRR-k-R#RC80sFRC#oH0RCs)7q7)H
#oDMNR8IN_osCR:RRR8#0_oDFHPO_CFO0s85N8HsI8-0E4FR8IFM0R;j2RRRRRR--k8#CRR0FsHCo#s0CR7Wq7#)
HNoMDFRDIN_s8R8s:0R#8F_Do_HOP0COFcs5RI8FMR0FjR2;RRRRRRRRRRRRR-R-R8sN8LsRHR0#HkMb0FR0Rv)qRDOCD5#R6HRL0s#RCHJks2C8
o#HMRNDD_FII8N8sRR:#_08DHFoOC_POs0F58cRF0IMF2Rj;RRRRRRRRRRRRRRR-I-RNs88R0LH#MRHbRk00)FRqOvRC#DDRR56L#H0RJsCkCHs802
$RbC0_lbNs88_b0$C#RHRsNsN5$RM_klODCD#C_8C8bRF0IMF2RjRRFV#_08DHFoOC_POs0FRR5g8MFI0jFR2#;
HNoMDlR0b8_N8RsR:lR0b8_N80s_$;bC
C
Lo
HM
RRRRR--QNVR8I8sHE80R6<RR#N#HRoM'Rj'0kFRMCk#8HRL0R#
RzRR4:RRRRHV58N8s8IH0=ERRR42oCCMsCN0
RRRRRRRRIDF_8sN8<sR=jR"j"jjRs&RNs8_Cjo52R;
RRRRRDRRFII_Ns88RR<="jjjj&"RR8IN_osC5;j2
RRRR8CMRMoCC0sNC4Rz;R
RR.RzRRR:H5VRNs88I0H8ERR=.o2RCsMCN
0CRRRRRRRRD_FIs8N8s=R<Rj"jj&"RR8sN_osC584RF0IMF2Rj;R
RRRRRRFRDIN_I8R8s<"=Rj"jjRI&RNs8_C4o5RI8FMR0Fj
2;RRRRCRM8oCCMsCN0R;z.
RRRRRzdRH:RVNR58I8sHE80Rd=R2CRoMNCs0RC
RRRRRDRRFsI_Ns88RR<=""jjRs&RNs8_C.o5RI8FMR0Fj
2;RRRRRRRRD_FII8N8s=R<Rj"j"RR&I_N8s5Co.FR8IFM0R;j2
RRRR8CMRMoCC0sNCdRz;R
RRcRzRRR:H5VRNs88I0H8ERR=co2RCsMCN
0CRRRRRRRRD_FIs8N8s=R<R''jRs&RNs8_Cdo5RI8FMR0Fj
2;RRRRRRRRD_FII8N8s=R<R''jRI&RNs8_Cdo5RI8FMR0Fj
2;RRRRCRM8oCCMsCN0R;zc
RRRRRz6RH:RVNR58I8sHE80Rc>R2CRoMNCs0RC
RRRRRDRRFsI_Ns88RR<=s_N8s5CocFR8IFM0R;j2
RRRRRRRRIDF_8IN8<sR=NRI8C_soR5c8MFI0jFR2R;
RCRRMo8RCsMCNR0Cz
6;
RRRRR--Q5VR8_HMs2CoRosCHC#0sQR7h#RkHRMoB
piRRRRzRnR:VRHRH58MC_soo2RCsMCN
0CRRRRRRRRbOsFCR##5iBp,QR7hL2RCMoH
RRRRRRRRRRRRRHV5iBpR'=R4N'RMB8RpCi'P0CM2ER0CRM
RRRRRRRRRRRRRHRRMC_so=R<Rj5"j"jjR7&RQ;h2
RRRRRRRRRRRR8CMR;HV
RRRRRRRR8CMRFbsO#C#;R
RRMRC8CRoMNCs0zCRnR;
RzRR(:RRRRHV50MFRM8H_osC2CRoMNCs0RC
RRRRRRRRRHRRMC_so=R<Rj5"j"jjR7&RQ;h2
RRRR8CMRMoCC0sNC(Rz;R

R-RR-VRQRN5s8_8ss2CoRosCHC#0sqR)7R7)kM#HopRBiR
RR4Rzj:RRRRHV58sN8ss_CRo2oCCMsCN0
RRRRRRRRFbsO#C#RB5mpRi,)7q7)L2RCMoH
RRRRRRRRRRRRRHV5pmBiRR='R4'NRM8miBp'CCPMR020MEC
RRRRRRRRRRRRRRRR8sN_osCRR<=)7q7)85N8HsI8-0E4FR8IFM0R;j2
RRRRRRRRRRRR8CMR;HV
RRRRRRRR8CMRFbsO#C#;R
RRMRC8CRoMNCs0zCR4
j;RRRRzR44:VRHRF5M0NRs8_8ss2CoRMoCC0sNCR
RRRRRRRRRRNRs8C_so=R<R7)q7N)58I8sHE80-84RF0IMF2Rj;R
RRMRC8CRoMNCs0zCR4
4;RRRRRRRR
RRRRR--Q5VRI8N8sC_sos2RC#oH0RCsW7q7)#RkHRMoB
piRRRRzR4.RH:RVIR5Ns88_osC2CRoMNCs0RC
RRRRRbRRsCFO#5#RB,piR7Wq7R)2LHCoMR
RRRRRRRRRRVRHRp5BiRR='R4'NRM8B'piCMPC002RE
CMRRRRRRRRRRRRRRRRI_N8sRCo<W=Rq)7758N8s8IH04E-RI8FMR0Fj
2;RRRRRRRRRRRRCRM8H
V;RRRRRRRRCRM8bOsFC;##
RRRR8CMRMoCC0sNC4Rz.R;
RzRR4:dRRRHV50MFR8IN8ss_CRo2oCCMsCN0
RRRRRRRRRRRR8IN_osCRR<=W7q7)R;
RCRRMo8RCsMCNR0Cz;4d
R
RR-R-RMtCC0sNCER0CqR)vCRODRD#NRM8#CCDOD0RFOoH
RRRRcz4RV:RFHsRRRHMM_klODCD#C_8C8bRF0IMFRRjoCCMsCN0
RRRRR--ADkH8kRF00bkRNCMLRDC#CCDOD0RFOoH
RRRRRRRRR--Q5VRNs88I0H8ERR>4R62O'NM0#RkCRRN1BpQRDOCDR
RRRRRR Rm4:nRRRHV58N8s8IH0>ERR246RMoCC0sNCR
RRRRRRRRRRRRRRkRF0M_C5RH2<'=R4I'RERCM58sN_osC58N8s8IH04E-RI8FMR0F6=2RRRH2CCD#R''j;R
RRRRRRMRC8CRoMNCs0mCR ;4n
RRRRRRRRR--Q5VRNs88I0H8ERR>6q2Rh57RNs88I0H8E=R<R246RNk#R1NRpRQBODCD
RRRRRRRR4m 6RR:H5VRNs88I0H8ERR=4R62oCCMsCN0
RRRRRRRRRRRRRRRRb0l_8N8s25H58gRF0IMF2RjRR<=h5maOPFM_8#0_oDFHPO_CFO0s,5HR24j2mRX)NRs8C_so85N8HsI8-0E4FR8IFM0R;62
RRRRRRRRRRRRRRRRh1q76_4R1:Rq4h7jFRbsl0RN5bRq>R=Rb0l_8N8s25H5,j2R=AR>lR0b8_N8Hs52254,RRB=0>RlNb_858sH.2527,RRR=>0_lbNs8855H2d
2,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR RRRR=>0_lbNs8855H2cR2,w>R=Rb0l_8N8s25H5,62R=tR>lR0b8_N8Hs5225n,RR]=0>RlNb_858sH(252
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRQRRRR=>0_lbNs8855H2UR2,K>R=Rb0l_8N8s25H5,g2R=ZR>kRF0M_C52H2;R
RRRRRRMRC8CRoMNCs0mCR ;46
RRRRRRRR4m cRR:H5VRNs88I0H8ERR=4Rc2oCCMsCN0
RRRRRRRRRRRRRRRRb0l_8N8s25H58URF0IMF2RjRR<=h5maOPFM_8#0_oDFHPO_CFO0s,5HR2g2R)XmR8sN_osC58N8s8IH04E-RI8FMR0F6
2;RRRRRRRRRRRRRRRR17qh_R4c:qR1hj74RsbF0NRlbqR5RR=>0_lbNs8855H2jR2,A>R=Rb0l_8N8s25H5,42R=BR>lR0b8_N8Hs5225.,RR7=0>RlNb_858sHd252R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR =0>RlNb_858sHc252w,RRR=>0_lbNs8855H26R2,t>R=Rb0l_8N8s25H5,n2R=]R>lR0b8_N8Hs5225(,RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRQ=0>RlNb_858sHU252K,RRR=>',4'R=ZR>kRF0M_C52H2;R
RRRRRRMRC8CRoMNCs0mCR ;4c
RRRRRRRR4m dRR:H5VRNs88I0H8ERR=4Rd2oCCMsCN0
RRRRRRRRRRRRRRRRb0l_8N8s25H58(RF0IMF2RjRR<=h5maOPFM_8#0_oDFHPO_CFO0s,5HR2U2R)XmR8sN_osC58N8s8IH04E-RI8FMR0F6
2;RRRRRRRRRRRRRRRR17qh_R4d:qR1hR7URsbF0NRlbqR5RR=>0_lbNs8855H2jR2,A>R=Rb0l_8N8s25H5,42R=BR>lR0b8_N8Hs5225.,RR7=0>RlNb_858sHd252R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR =0>RlNb_858sHc252w,RRR=>0_lbNs8855H26R2,t>R=Rb0l_8N8s25H5,n2R=]R>lR0b8_N8Hs5225(,RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRZ=F>RkC0_M25H2R;
RRRRRCRRMo8RCsMCNR0Cmd 4;R
RRRRRR Rm4:.RRRHV58N8s8IH0=ERR24.RMoCC0sNCR
RRRRRRRRRRRRRRlR0b8_N8Hs52R5n8MFI0jFR2=R<Rahm5MOFP0_#8F_Do_HOP0COFHs5,2R(2mRX)NRs8C_so85N8HsI8-0E4FR8IFM0R;62
RRRRRRRRRRRRRRRRh1q7._4R1:RqUh7RFRbsl0RN5bRq>R=Rb0l_8N8s25H5,j2R=AR>lR0b8_N8Hs52254,RRB=0>RlNb_858sH.2527,RRR=>0_lbNs8855H2d
2,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR RRRR=>0_lbNs8855H2cR2,w>R=Rb0l_8N8s25H5,62R=tR>lR0b8_N8Hs5225n,RR]='>R4R',
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRZ>R=R0Fk_5CMH;22
RRRRRRRR8CMRMoCC0sNC Rm4
.;RRRRRRRRm4 4RH:RVNR58I8sHE80R4=R4o2RCsMCN
0CRRRRRRRRRRRRRRRR0_lbNs8855H26FR8IFM0RRj2<h=RmOa5F_MP#_08DHFoOC_POs0F5RH,nR22XRm)s_N8s5CoNs88I0H8ER-48MFI06FR2R;
RRRRRRRRRRRRR1RRq_h74:4RRh1q7RnRb0FsRblNRR5q=0>RlNb_858sHj252A,RRR=>0_lbNs8855H24R2,B>R=Rb0l_8N8s25H5,.2R=7R>lR0b8_N8Hs5225d,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR= R>lR0b8_N8Hs5225c,RRw=0>RlNb_858sH6252Z,RRR=>F_k0CHM52
2;RRRRRRRRCRM8oCCMsCN0R4m 4R;
RRRRRmRR R4j:VRHR85N8HsI8R0E=jR42CRoMNCs0RC
RRRRRRRRRRRRR0RRlNb_858sHc25RI8FMR0Fj<2R=mRhaF5OM#P_0D8_FOoH_OPC05FsH6,R2X2Rms)RNs8_CNo58I8sHE80-84RF0IMF2R6;R
RRRRRRRRRRRRRRqR1h47_jRR:17qhnbRRFRs0lRNb5=qR>lR0b8_N8Hs5225j,RRA=0>RlNb_858sH4252B,RRR=>0_lbNs8855H2.R2,7>R=Rb0l_8N8s25H5,d2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR >R=Rb0l_8N8s25H5,c2R=wR>4R''Z,RRR=>F_k0CHM52
2;RRRRRRRRCRM8oCCMsCN0R4m jR;
RRRRRmRR RgR:VRHR85N8HsI8R0E=2RgRMoCC0sNCR
RRRRRRRRRRRRRRlR0b8_N8Hs52R5d8MFI0jFR2=R<Rahm5MOFP0_#8F_Do_HOP0COFHs5,2Rc2mRX)NRs8C_so85N8HsI8-0E4FR8IFM0R;62
RRRRRRRRRRRRRRRRh1q7R_g:qR1hR7cRFRbsl0RN5bRq>R=Rb0l_8N8s25H5,j2R=AR>lR0b8_N8Hs52254,RRB=0>RlNb_858sH.2527,RRR=>0_lbNs8855H2d
2,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRZRRRR=>F_k0CHM52
2;RRRRRRRRCRM8oCCMsCN0Rgm ;R
RRRRRR RmU:RRRRHV58N8s8IH0=ERRRU2oCCMsCN0
RRRRRRRRRRRRRRRRb0l_8N8s25H58.RF0IMF2RjRR<=h5maOPFM_8#0_oDFHPO_CFO0s,5HR2d2R)XmR8sN_osC58N8s8IH04E-RI8FMR0F6
2;RRRRRRRRRRRRRRRR17qh_:URRh1q7RcRRsbF0NRlbqR5RR=>0_lbNs8855H2jR2,A>R=Rb0l_8N8s25H5,42R=BR>lR0b8_N8Hs5225.,RR7='>R4
',RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRZRRRR=>F_k0CHM52
2;RRRRRRRRCRM8oCCMsCN0RUm ;R
RRRRRR Rm(:RRRRHV58N8s8IH0=ERRR(2oCCMsCN0
RRRRRRRRRRRRRRRRb0l_8N8s25H584RF0IMF2RjRR<=h5maOPFM_8#0_oDFHPO_CFO0s,5HR2.2R)XmR8sN_osC58N8s8IH04E-RI8FMR0F6
2;RRRRRRRRRRRRRRRR17qh_:(RRh1q7R.RRsbF0NRlbqR5RR=>0_lbNs8855H2jR2,A>R=Rb0l_8N8s25H5,42R=ZR>kRF0M_C52H2;R
RRRRRRMRC8CRoMNCs0mCR 
(;RRRRRRRRmR nRH:RVNR58I8sHE80Rn=R2CRoMNCs0RC
RRRRRRRRRRRRRFRRkC0_M25HRR<='R4'IMECRN5s8C_so256RO=RF_MP#_08DHFoOC_POs0F54H,225j2DRC#'CRj
';RRRRRRRRCRM8oCCMsCN0Rnm ;R
RR-R-RRQV58N8s8IH0<ER=2R6RRMFFbk0kC0RMDNLCCR#D0CORoDFHMORCCC88R
RRRRRR Rm6RR:H5VRNs88I0H8E=R<RR62oCCMsCN0
RRRRRRRRRRRRRRRR0Fk_5CMH<2R=4R''R;
RRRRRCRRMo8RCsMCNR0Cm; 6
R
RR-R-RRQV58N8s8IH0>ERRRg2kR#CWju RR0F8FCO8NCR8C8s#L#RHR0#nER0soFkERRgNRM8W4u RR0F8FCO8LCRHR0#4+jR
RRRRRRRR4W jRR:H5VRNs88I0H8ERR>go2RCsMCN
0CRRRRRRRRRRRRRRRRIjbC_5CMH<2R=4R''ERIC5MRI_N8s5CoUFR8IFM0RR62=FROM#P_0D8_FOoH_OPC05FsHj,.2R5d8MFI0jFR2C2RDR#C';j'
RRRRRRRRRRRRRRRRCIb4M_C5RH2<'=R4I'RERCM58IN_osC58N8s8IH04E-RI8FMR0Fg=2RRMOFP0_#8F_Do_HOP0COFHs5,2.j58N8s8IH0nE-RI8FMR0FcR22CCD#R''j;R
RRRRRRRRRRMRC8CRoMNCs0WCR ;4j
RRRRR--Q5VRNs88I0H8ERR=UsRFRRg2kR#CWju RR0F8FCO8NCR8C8s#L#RHR0#nER0soFkE
RgRRRRRRRRWR gRH:RV5R5Ns88I0H8ERR=Um2R)NR58I8sHE80Rg=R2o2RCsMCN
0CRRRRRRRRRRRRRRRRIjbC_5CMH<2R=4R''ERIC5MRI_N8s5CoNs88I0H8ER-48MFI06FR2RR=HC2RDR#C';j'
RRRRRRRRRRRRRRRRCIb4M_C5RH2<'=R4
';RRRRRRRRRRRRCRM8oCCMsCN0RgW ;R
RR-R-RRQV58N8s8IH0=ERRR(2kR#CWju RR0F8FCO80CREnCR0NER8C8s#L#RH&0RR Wu4FR0RO8CFR8C0REC(R0ENs88CR##L
H0RRRRRRRRWR (RH:RVNR58I8sHE80R(=R2CRoMNCs0RC
RRRRRRRRRRRRRIRRb_CjCHM52=R<R''4RCIEMIR5Ns8_C6o52RR=OPFM_8#0_oDFHPO_CFO0s,5H.j252C2RDR#C';j'
RRRRRRRRRRRRRRRRCIb4M_C5RH2<'=R4I'RERCM58IN_osC5Rn2=FROM#P_0D8_FOoH_OPC05FsH2,.5242R#CDCjR''R;
RRRRRCRRMo8RCsMCNR0CW; (
RRRRR--Q5VRNs88I0H8ERR=nk2R#WCRuR j08FRC8OFCER0C0RnE8RN8#sC#HRL0R
RRRRRR RWn:RRRRHV58N8s8IH0=ERRRn2oCCMsCN0
RRRRRRRRRRRRRRRRCIbjM_C5RH2<'=R4I'RERCM58IN_osC5R62=FROM#P_0D8_FOoH_OPC05FsH2,452j2R#CDCjR''R;
RRRRRRRRRRRRRIRRb_C4CHM52=R<R''4;R
RRRRRRMRC8CRoMNCs0WCR 
n;RRRR-Q-RVNR58I8sHE80RR<=6M2RFsRIHR0CCLMND#CRCODC0FRDoRHOM8CCCR8
RRRRRWRR R6R:VRHR85N8HsI8R0E<6=R2CRoMNCs0RC
RRRRRRRRRRRRRIRRb_CjCHM52=R<R''4;R
RRRRRRRRRRRRRRbRICC4_M25HRR<=';4'
RRRRRRRR8CMRMoCC0sNC RW6
;
RRRRCRM8oCCMsCN0Rcz4;R

RbRRsCFO#5#RB,piRh7Q2CRLo
HMRRRRRHRRVBR5p=iRR''4R8NMRiBp'CCPMR020MEC
RRRRRRRRRRRHsM_CRo4<H=RMC_soR;
RRRRRRRRR RW_t) 4=R<R;W 
RRRRRRRCRM8H
V;RRRRCRM8bOsFC;##
R
RR.Rz6RR:H5VRMRF080Fk_osC2CRoMNCs0RC
RRRRRzRR4:(4RFbsO#C#R 5W_t) 4),Rq)77,qRW7,7)R_HMs4Co,kRF0C_soR2
RRRRRLRRCMoH
RRRRRRRRRRRRRHV5 5W_t) 4RR='24'R8NMRq5)7R7)=qRW727)2ER0CRM
RRRRRRRRRRRRR7RRmRza<H=RMC_soI45HE80-84RF0IMF2Rj;R
RRRRRRRRRRDRC#RC
RRRRRRRRRRRRR7RRmRza<F=Rks0_CIo5HE80-84RF0IMF2Rj;R
RRRRRRRRRRMRC8VRH;R
RRRRRRMRC8sRbF#OC#4Rz(
4;RRRRCRM8oCCMsCN0R6z.;R

RzRRdRjR:VRHRF58ks0_CRo2oCCMsCN0
RRRRRRRRFbsO#C#RB5mpRi,F_k0s2CoRoLCHRM
RRRRRRRRRHRRVmR5BRpi=4R''MRN8BRmpCi'P0CM2ER0CRM
RRRRRRRRRRRRR7RRmRza<F=Rks0_CIo5HE80-84RF0IMF2Rj;R
RRRRRRRRRRMRC8VRH;R
RRRRRRMRC8sRbF#OC#R;
RCRRMo8RCsMCNR0Cz;dj
R
RR-R-RCtMsCN0RC0ERv)qRDOCDI#RHR0E0-sH#00NCR#
RzRR4:6RRsVFRHHRMkRMlC_OD_D#8bCCRI8FMR0FjCRoMNCs0RC
RRRRRzRR4:(RRsVFRH[RMkRMlC_OD_D#ICH8RI8FMR0FjCRoMNCs0RC
RRRRRRRRRzRR):qvR 7Bdc.XRR
RRRRRRRRRRRRRRFRbsl0RN5bR7RQj=H>RMC_so[55*2c2,QR74>R=R_HMs5Co5c[*22+4,QR7.>R=R_HMs5Co5c[*22+.,QR7d>R=R_HMs5Co5c[*22+d,R
RRRRRRRRRRRRRRRRRRRRRRRRRWjq7RR=>D_FII8N8s25j,qRW7=4R>FRDIN_I858s4R2,W.q7RR=>D_FII8N8s25.,qRW7=dR>FRDIN_I858sdR2,Wcq7RR=>D_FII8N8s25c,R
RRRRRRRRRRRRRRRRRRRRRRRRR)jq7RR=>D_FIs8N8s25j,qR)7=4R>FRDIN_s858s4R2,).q7RR=>D_FIs8N8s25.,qR)7=dR>FRDIN_s858sdR2,)cq7RR=>D_FIs8N8s25c,-
-RRRRRRRRRRRRRRRRRRRRRRRRR)RW =hR> RW,uRW =jR>bRICCj_M25H,uRW =4R>bRICC4_M25H,iRBRR=>h5maB2pi,RR
RRRRRRRRRRRRRRRRRRRRRRRRR W)h>R=R,W R Wuj>R=RCIbjM_C5,H2R Wu4>R=RCIb4M_C5,H2RRBi=B>RpRi,
RRRRRRRRRRRRRRRRRRRRRRRR7RRm=jR>kRF0k_L#,5H5c[*2R2,7Rm4=F>RkL0_kH#5,*5[c42+27,Rm=.R>kRF0k_L#,5H5c[*22+.,mR7d>R=R0Fk_#Lk55H,[2*c+2d2;R
RRRRRRRRRRRRRRkRF0C_so[55*2c2RR<=F_k0L5k#H[,5*2c2RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_so[55*+c24<2R=kRF0k_L#,5H5c[*22+4RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_so[55*+c2.<2R=kRF0k_L#,5H5c[*22+.RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_so[55*+c2d<2R=kRF0k_L#,5H5c[*22+dRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRMRC8CRoMNCs0zCR4
(;RRRRCRM8oCCMsCN0R6z4;-

-zRR.:URRRHV5k8F0C_soo2RCsMCN
0C-R-RRRRRR4RznRR:VRFsHMRHRlMk_DOCD8#_CRCb8MFI0jFRRMoCC0sNC-
-RRRRRRRRzR4U:FRVsRR[HMMRkOl_C#DD_8IHCFR8IFM0RojRCsMCN
0C-R-RRRRRRRRRR)RzqRv:7dB .RXc
R--RRRRRRRRRRRRRbRRFRs0lRNb5j7QRR=>HsM_C5o5[2*c27,RQ=4R>MRH_osC5*5[c42+27,RQ=.R>MRH_osC5*5[c.2+27,RQ=dR>MRH_osC5*5[cd2+2-,
-RRRRRRRRRRRRRRRRRRRRRRRRWRRqR7j=D>RFII_Ns885,j2R7Wq4>R=RIDF_8IN84s52W,RqR7.=D>RFII_Ns885,.2R7Wqd>R=RIDF_8IN8ds52W,RqR7c=D>RFII_Ns885,c2
R--RRRRRRRRRRRRRRRRRRRRRRRRR7)qj>R=RIDF_8sN8js52),RqR74=D>RFsI_Ns885,42R7)q.>R=RIDF_8sN8.s52),RqR7d=D>RFsI_Ns885,d2R7)qc>R=RIDF_8sN8cs52-,
-RRRRRRRRRRRRRRRRRRRRRRRRWRR)R h=W>R W,RuR j=I>Rb_CjCHM52W,RuR 4=I>Rb_C4CHM52B,Ri>R=Rahm5iBp2
,R-R-RRRRRRRRRRRRRRRRRRRRRRRRRTj7mRR=>F_k0L5k#H[,5*2c2,7RTm=4R>kRF0k_L#,5H5c[*22+4,7RTm=.R>kRF0k_L#,5H5c[*22+.,7RTm=dR>kRF0k_L#,5H5c[*22+d2-;
--
-RRRRRRRRRRRRRkRF0C_so[55*2c2RR<=F_k0L5k#H[,5*2c2RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;-
-RRRRRRRRRRRRRRRRF_k0s5Co5c[*22+4RR<=F_k0L5k#H[,5*+c24I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';-R-RRRRRRRRRRRRRRkRF0C_so[55*+c2.<2R=kRF0k_L#,5H5c[*22+.RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;-
-RRRRRRRRRRRRRRRRF_k0s5Co5c[*22+dRR<=F_k0L5k#H[,5*+c2dI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';-R-RRRRRRRRRRMRC8CRoMNCs0zCR4
U;-R-RRRRRR8CMRMoCC0sNC4Rzn-;
-RRRR8CMRMoCC0sNC.RzU
;
-R-RRRRRk:URRRHV5k8F0C_soo2RCsMCN
0C-R-RRRRR7amzRR<=F_k0s5CoI0H8ER-48MFI0jFR2-;
-CRRMo8RCsMCNR0Ck
U;RRRRRRRR
8CMRONsECH0Os0kCsRNO;Ej




