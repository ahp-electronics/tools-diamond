library verilog;
use verilog.vl_types.all;
entity config_jtag is
    port(
        prog_128        : in     vl_logic;
        idcode          : in     vl_logic_vector(31 downto 0);
        clear_finish    : in     vl_logic;
        por             : in     vl_logic;
        tms             : in     vl_logic;
        tck             : in     vl_logic;
        tdi             : in     vl_logic;
        asrout_0        : in     vl_logic;
        dsrout_0        : in     vl_logic;
        bsout_0         : in     vl_logic;
        cmd_ld_ucode    : in     vl_logic;
        cmd_prgm_done_r : in     vl_logic;
        cmd_prgm_done_comp: in     vl_logic;
        cmd_prgm_sec    : in     vl_logic;
        cmd_ld_ctrl0    : in     vl_logic;
        crc_err         : in     vl_logic;
        id_fail_r       : in     vl_logic;
        program         : in     vl_logic;
        mux_clk         : in     vl_logic;
        wakeup_clk      : in     vl_logic;
        cmd_ctrl0_r     : in     vl_logic_vector(31 downto 0);
        cmd_ucode_r     : in     vl_logic_vector(31 downto 0);
        er1out          : in     vl_logic;
        er2out          : in     vl_logic;
        clear_memory    : in     vl_logic;
        pll_lock        : in     vl_logic_vector(3 downto 0);
        ext_done        : in     vl_logic;
        forcearch_cfg   : in     vl_logic;
        done_phase      : in     vl_logic_vector(3 downto 0);
        goe_phase       : in     vl_logic_vector(2 downto 0);
        gwd_phase       : in     vl_logic_vector(2 downto 0);
        gsr_phase       : in     vl_logic_vector(2 downto 0);
        pll_set         : in     vl_logic_vector(3 downto 0);
        flash_status    : in     vl_logic;
        flash_fail      : in     vl_logic;
        syn_ext_done    : in     vl_logic;
        toe             : in     vl_logic;
        all_dwnld_done  : in     vl_logic;
        cfg             : in     vl_logic_vector(1 downto 0);
        wakeup          : out    vl_logic;
        mclk_en_r       : out    vl_logic;
        jtag_state      : out    vl_logic_vector(3 downto 0);
        jtag_active     : out    vl_logic;
        edit_mod        : out    vl_logic;
        auto_clear_en   : out    vl_logic;
        mck_freq_switch : out    vl_logic;
        jtag_data       : out    vl_logic;
        jtag_addr       : out    vl_logic;
        tdo_out         : out    vl_logic;
        tdo_en          : out    vl_logic;
        done_pupb       : out    vl_logic;
        freq_sel        : out    vl_logic_vector(5 downto 0);
        freq_div        : out    vl_logic_vector(5 downto 0);
        init_r          : out    vl_logic;
        rst_addr_o      : out    vl_logic;
        rti             : out    vl_logic;
        goe_high_r      : out    vl_logic;
        gwd_high_r      : out    vl_logic;
        gsr_high_r      : out    vl_logic;
        done_high_all   : out    vl_logic;
        selasr          : out    vl_logic;
        seldsr          : out    vl_logic;
        read_o          : out    vl_logic;
        vfy_incr_rti_o  : out    vl_logic;
        bsmode1         : out    vl_logic;
        bsmode2         : out    vl_logic;
        bsmode3         : out    vl_logic;
        wakeup_minus_r  : out    vl_logic;
        wakeup_minus    : out    vl_logic;
        jtag_unprogram  : out    vl_logic;
        jtag_functional : out    vl_logic;
        shiftdr         : out    vl_logic;
        upir            : out    vl_logic;
        capdr           : out    vl_logic;
        updr            : out    vl_logic;
        seldr           : out    vl_logic;
        selir           : out    vl_logic;
        tlreset         : out    vl_logic;
        done_reg        : out    vl_logic;
        extest          : out    vl_logic;
        sample          : out    vl_logic;
        selbsr          : out    vl_logic;
        mfg_bits        : out    vl_logic_vector(179 downto 0);
        init            : out    vl_logic;
        refresh_o       : out    vl_logic;
        erase_ee_o      : out    vl_logic;
        erase_sram_o    : out    vl_logic;
        eraseall_ee_o   : out    vl_logic;
        eraseall_sram_o : out    vl_logic;
        ucode_ee_o      : out    vl_logic;
        edit_tran       : out    vl_logic;
        program_ee_o    : out    vl_logic;
        program_sram_o  : out    vl_logic;
        prog_inc_rti_ee_o: out    vl_logic;
        prog_inc_rti_sram_o: out    vl_logic;
        progucode_ee_o  : out    vl_logic;
        progpes_ee_o    : out    vl_logic;
        progsec_ee_o    : out    vl_logic;
        progdone_ee_o   : out    vl_logic;
        read_pes_o      : out    vl_logic;
        vfy_incr_rti_ee_o: out    vl_logic;
        read_ee_o       : out    vl_logic;
        ee_mod          : out    vl_logic;
        fl_edit_dwnld   : out    vl_logic;
        program_effect  : out    vl_logic;
        j_fl_ep         : out    vl_logic;
        mfg_prg_red     : out    vl_logic;
        read_dnld_red   : out    vl_logic;
        verify_jtag     : out    vl_logic;
        j_fl_ep_only    : out    vl_logic;
        mc1_goe_en      : in     vl_logic;
        usr_goe         : in     vl_logic;
        erase_tag_o     : out    vl_logic;
        prog_tag_o      : out    vl_logic;
        read_tag_o      : out    vl_logic;
        e2_secty        : out    vl_logic;
        ues_crc_dsr     : out    vl_logic_vector(31 downto 0);
        erase_pulse     : in     vl_logic;
        flash_mini      : in     vl_logic_vector(205 downto 0);
        flash_sec_l     : in     vl_logic_vector(3 downto 0);
        latch_encr      : in     vl_logic;
        latch_shadow    : in     vl_logic;
        done_ee_r       : out    vl_logic;
        mfg_era_red     : out    vl_logic;
        jtag_store      : out    vl_logic;
        cfg_dd          : in     vl_logic;
        program_spi     : out    vl_logic;
        chip_crc_2_reg  : in     vl_logic_vector(31 downto 0);
        cmd_st_crc32    : in     vl_logic;
        sed_rdbk        : in     vl_logic;
        spisi           : in     vl_logic;
        ssi_en          : in     vl_logic;
        sso_en          : in     vl_logic;
        chip_crc_fm_reg : out    vl_logic_vector(31 downto 0);
        sso             : out    vl_logic;
        progcrc32_ee_o  : out    vl_logic;
        read_crc_ee_o   : out    vl_logic;
        sspi_capdr      : in     vl_logic;
        sspi_idcode_o   : in     vl_logic;
        sspi_progcrc32_ee_o: in     vl_logic;
        sspi_progctrl0_ee_o: in     vl_logic;
        sspi_progucode_ee_o: in     vl_logic;
        sspi_ucode_ee_o : in     vl_logic;
        sspi_ucode_o    : in     vl_logic;
        sspi_vfycrc32_ee_o: in     vl_logic;
        sspi_vfycrc32_o : in     vl_logic;
        sspi_vfyctrl0_ee_o: in     vl_logic;
        sspi_vfyctrl0_o : in     vl_logic;
        spi_prgm_clear  : out    vl_logic;
        async_rst       : out    vl_logic;
        prem_time_out   : in     vl_logic;
        sed_enable_nedge: in     vl_logic;
        nonjtag_cfg_r   : in     vl_logic;
        sospi           : in     vl_logic;
        freeze_io_en    : out    vl_logic;
        auto_rconf      : in     vl_logic;
        status_out      : in     vl_logic;
        status_cap      : out    vl_logic;
        status_shift    : out    vl_logic;
        decrypt_o       : out    vl_logic;
        erase_encr_ee_o : out    vl_logic;
        prog_encr_ee_o  : out    vl_logic;
        read_encr_ee_o  : out    vl_logic;
        encrypt_r       : out    vl_logic_vector(127 downto 0);
        otp_active      : out    vl_logic;
        sspi_refresh_o  : in     vl_logic;
        shf128_r        : out    vl_logic_vector(127 downto 0);
        decrypt_en      : out    vl_logic;
        sspi_decrypt_o  : in     vl_logic;
        sspi_protect_o  : in     vl_logic;
        sf_secty        : out    vl_logic;
        dsrout_tag      : in     vl_logic;
        sspi_progsec_ee_o: in     vl_logic;
        sspi_read_tag_o : in     vl_logic;
        sed_prgm_n      : in     vl_logic;
        key_r           : out    vl_logic;
        reset_crc16     : out    vl_logic;
        cmd_crc         : in     vl_logic_vector(15 downto 0);
        sspi_rdstatus   : in     vl_logic;
        sspi_read_crc16 : in     vl_logic;
        cap_bp          : out    vl_logic;
        seler1          : out    vl_logic;
        seler2          : out    vl_logic;
        sspi_progdis_o  : in     vl_logic;
        edit_tran_cdu   : out    vl_logic;
        flclk           : in     vl_logic
    );
end config_jtag;
