library verilog;
use verilog.vl_types.all;
entity HCLK_TREE is
    port(
        A               : in     vl_logic;
        Z               : out    vl_logic
    );
end HCLK_TREE;
