--
@ER--B$FbsEHo0OR52gR4g-cRRj.jd$R1MHbDO$H0ROQM
R--fN]C8:CsR#//$DMbH0OH$N/lb..jjDjdNl0/NCbbsN#/0D0/HoL/CFM_scONCN/slI_s38PEyf4R

--
-
-

---1-RHDlbCqR)vHRI0#ERHDMoC7Rq71) 1FRVsCRsNN8RMI8RsCH0
R--aoNsC:0RROpkCRM0-)RmBcqR -
-
LDHs$NsRCHCCk;
#HCRC3CC#_08DHFoO4_4nNc3D
D;kR#CHCCC38#0_oDFH#O_HCoM8D3NDk;
#HCRC3CC#_08DHFoOs_NH30EN;DD
D--HNLssF$RscON;-
-kR#CFNsOcs3FOFNOlNb3D
D;-0-N0LsHkR0C#_$MLODN	F_LGVRFR )Bdc.XRO:RFFlbM0CMRRH#0Csk;C

M00H$qR)vW_)R
H#RRRRoCCMsRHO5R
RRRRRRNRVl$HD:0R#soHMRR:="MMFC
";RRRRRRRRI0H8ERR:HCM0oRCs:(=R;RR
RRRRRNRR8I8sHE80RH:RMo0CC:sR=;R(RRRRRRRR-L-RHCoRMoFkEFRVsCR8b
0ERRRRRRRR80CbERR:HCM0oRCs:R=R4;.U
RRRRRRRRk8F0C_soRR:LDFFCRNM:V=RNCD#;RRRR-R-R#ENR0FkbRk0s
CoRRRRRRRR8_HMsRCo:FRLFNDCM=R:RDVN#RC;RRRRRR--ERN#8NN0RbHMks0RCRo
RRRRRNRR8_8ssRCo:FRLFNDCM=R:RDVN#RCRRRRR-E-RNs8RCRN8Ns88CR##s
CoRRRRRRRR2R;
RbRRFRs05R
RRRRRRmR7zRaR:kRF00R#8F_Do_HOP0COFIs5HE80-84RF0IMF2Rj;R
RRRRRRQR7hRRR:MRHR0R#8F_Do_HOP0COFIs5HE80-84RF0IMF2Rj;R
RRRRRR7Rq7R)R:MRHR0R#8F_Do_HOP0COFNs58I8sHE80-84RF0IMF2Rj;R
RRRRRR RWRRRR:MRHR0R#8F_Do;HORRRRR-RR-sRIHR0CCLMNDVCRFssRNRl
RRRRRBRRpRiRRH:RM#RR0D8_FOoH;RRRRRRR-O-RD	FORsVFRlsN,8RN8Rs,8
HMRRRRRRRRmiBpRRR:HRMR#_08DHFoORRRRRRRRR--FRb0OODF	FRVsFR8kR0
RRRRR2RR;M
C8MRC0$H0Rv)q_;)W
-
-
R--w#Hs0lRHblDCCNM00MHFR#lk0CRLRDONDRC8NEsOj-
-
ONsECH0Os0kCsRNOREjF)VRq)v_W#RH
lOFbCFMM10RqUh7
FRbs50R
RRRqRR:H#MR0D8_FOoH;R
RR:ARRRHM#_08DHFoOR;
RRRB:MRHR8#0_oDFH
O;R7RRRH:RM0R#8F_Do;HO
RRR RR:H#MR0D8_FOoH;R
RR:wRRRHM#_08DHFoOR;
RRRt:MRHR8#0_oDFH
O;R]RRRH:RM0R#8F_Do;HO
RRRZRR:FRk0#_08DHFoO2
R;M
C8FROlMbFC;M0
lOFbCFMM10Rqnh7
FRbs50R
RRRqRR:H#MR0D8_FOoH;R
RR:ARRRHM#_08DHFoOR;
RRRB:MRHR8#0_oDFH
O;R7RRRH:RM0R#8F_Do;HO
RRR RR:H#MR0D8_FOoH;R
RR:wRRRHM#_08DHFoOR;
RRRZ:kRF00R#8F_Do
HOR
2;CRM8ObFlFMMC0O;
FFlbM0CMRh1q7Rc
b0FsRR5
RRRq:MRHR8#0_oDFH
O;RARRRH:RM0R#8F_Do;HO
RRRBRR:H#MR0D8_FOoH;R
RR:7RRRHM#_08DHFoOR;
RRRZ:kRF00R#8F_Do
HOR
2;CRM8ObFlFMMC0O;
FFlbM0CMRh1q7R.
b0FsRR5
RRRq:MRHR8#0_oDFH
O;RARRRH:RM0R#8F_Do;HO
RRRZRR:FRk0#_08DHFoO2
R;M
C8FROlMbFC;M0
F
OlMbFCRM017qh4Rj
b0FsRR5
RRRq:MRHR8#0_oDFH
O;RARRRH:RM0R#8F_Do;HO
RRRBRR:H#MR0D8_FOoH;R
RR:7RRRHM#_08DHFoOR;
RRR :MRHR8#0_oDFH
O;RwRRRH:RM0R#8F_Do;HO
RRRtRR:H#MR0D8_FOoH;R
RR:]RRRHM#_08DHFoOR;
RRRQ:MRHR8#0_oDFH
O;RKRRRH:RM0R#8F_Do;HO
RRRZRR:FRk0#_08DHFoO2
R;M
C8FROlMbFC;M0
lOFbCFMM)0RB. dXRc
b0FsRR5
R7RqjRR:H#MR0D8_FOoH;R
RR4q7RH:RM0R#8F_Do;HO
RRRqR7.:MRHR8#0_oDFH
O;RqRR7:dRRRHM#_08DHFoOR;
R7RqcRR:H#MR0D8_FOoH;R
RRj7QRH:RM0R#8F_Do;HO
RRR7RQ4:MRHR8#0_oDFH
O;R7RRQ:.RRRHM#_08DHFoOR;
RQR7dRR:H#MR0D8_FOoH;R
RRRBi:MRHR8#0_oDFH
O;RtRR1:)RRRHM#_08DHFoOR;
R)RW :hRRRHM#_08DHFoOR;
RuRW :jRRRHM#_08DHFoOR;
RuRW :4RRRHM#_08DHFoOR;
RmR7jRR:FRk0#_08DHFoOR;
RmR74RR:FRk0#_08DHFoOR;
RmR7.RR:FRk0#_08DHFoOR;
RmR7dRR:FRk0#_08DHFoOR;
R7RTm:jRR0FkR8#0_oDFH
O;RTRR7Rm4:kRF00R#8F_Do;HO
RRRT.7mRF:Rk#0R0D8_FOoH;R
RRmT7dRR:FRk0#_08DHFoO2
R;M
C8FROlMbFC;M0
MOF#M0N0kRMlC_OD_D#8bCCRH:RMo0CC:sR=5R580CbERR-4d2/.R2;RRRRRRRR-y-RRRFVs#FIRRFV)dB .RXcODCD#CRMC88C
MOF#M0N0kRMlC_OD_D#ICH8RH:RMo0CC:sR=5R5I0H8ERR-4c2/2R;RRRRRRRRR-y-RRRFVOkFDlRM#F)VRB. dXOcRC#DDRCMC8
C80C$bR0Fk_#Lk_b0$C#RHRsNsN5$RM_klODCD#C_8C8bRF0IMF,RjRk5MlC_OD_D#ICH8*+c2dFR8IFM0RRj2F#VR0D8_FOoH;H
#oDMNR0Fk_#LkR:RRR0Fk_#Lk_b0$CR;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--.N7Rs$sNRRFV80FkRM5HbRk000FRs#H-0CN0##2
HNoMDkRF0M_CRRRR:0R#8F_Do_HOP0COFMs5kOl_C#DD_C8CbFR8IFM0R;j2R-R-RNCML#DCRsVFRH0s-N#00
C##MHoNIDRb_CjCRMRR#:R0D8_FOoH_OPC05FsM_klODCD#C_8C8bRF0IMF2Rj;-RR-sRIHR0CCLMNDRC#VRFsCENORIsFRRFV)RqvODCD#H
#oDMNRCIb4M_CR:RRR8#0_oDFHPO_CFO0sk5MlC_OD_D#8bCCRI8FMR0FjR2;RR--I0sHCMRCNCLD#FRVsNRCOsERFFIRVqR)vCROD
D##MHoNHDRMC_soRRRR#:R0D8_FOoH_OPC05FsI0H8ER+d8MFI0jFR2R;RRRRRR-RR-#RkC08RFCRso0H#C7sRQ
hR#MHoNFDRks0_CRoRR#:R0D8_FOoH_OPC05FsI0H8ER+d8MFI0jFR2R;RRRRRR-RR-#RkC08RFCRso0H#C7sRm
za#MHoNHDRMC_soR4RR#:R0D8_FOoH_OPC05FsI0H8ER+d8MFI0jFR2R;RR#R
HNoMD8RN_osCRRRR:0R#8F_Do_HOP0COFNs58I8sHE80-84RF0IMF2Rj;RRRR-R-RCk#8FR0RosCHC#0s7Rq7#)
HNoMDFRDI8_N8RsR:0R#8F_Do_HOP0COFcs5RI8FMR0FjR2;RRRRRRRRRRRRR-R-R8N8sHRL0H#RM0bkRR0F)RqvODCD#6R5R0LH#CRsJskHC
820C$bRb0l_8N8s$_0bHCR#sRNsRN$5lMk_DOCD8#_CRCb8MFI0jFR2VRFR8#0_oDFHPO_CFO0sgR5RI8FMR0Fj
2;#MHoN0DRlNb_8R8sR0:RlNb_8_8s0C$b;L

CMoH
R
RR-R-RRQVNs88I0H8ERR<6#RN#MHoR''jRR0Fk#MkCL8RH
0#RRRRzR4R:VRHR85N8HsI8R0E=2R4RMoCC0sNCR
RRRRRRFRDI8_N8<sR=jR"j"jjRN&R8C_so25j;R
RRMRC8CRoMNCs0zCR4R;
RzRR.:RRRRHV58N8s8IH0=ERRR.2oCCMsCN0
RRRRRRRRIDF_8N8s=R<Rj"jj&"RR_N8s5Co4FR8IFM0R;j2
RRRR8CMRMoCC0sNC.Rz;R
RRdRzRRR:H5VRNs88I0H8ERR=do2RCsMCN
0CRRRRRRRRD_FINs88RR<=""jjRN&R8C_soR5.8MFI0jFR2R;
RCRRMo8RCsMCNR0Cz
d;RRRRzRcR:VRHR85N8HsI8R0E=2RcRMoCC0sNCR
RRRRRRFRDI8_N8<sR=jR''RR&Ns8_Cdo5RI8FMR0Fj
2;RRRRCRM8oCCMsCN0R;zc
RRRRRz6RH:RVNR58I8sHE80Rc>R2CRoMNCs0RC
RRRRRDRRFNI_8R8s<N=R8C_soR5c8MFI0jFR2R;
RCRRMo8RCsMCNR0Cz
6;
RRRRR--Q5VR8_HMs2CoRosCHC#0sQR7h#RkHRMoB
piRRRRzRnR:VRHRH58MC_soo2RCsMCN
0CRRRRRRRRbOsFCR##5iBp,QR7hL2RCMoH
RRRRRRRRRRRRRHV5iBpR'=R4N'RMB8RpCi'P0CM2ER0CRM
RRRRRRRRRRRRRHRRMC_so=R<Rj5"j"jjR7&RQ;h2
RRRRRRRRRRRR8CMR;HV
RRRRRRRR8CMRFbsO#C#;R
RRMRC8CRoMNCs0zCRnR;
RzRR(:RRRRHV50MFRM8H_osC2CRoMNCs0RC
RRRRRRRRRHRRMC_so=R<Rj5"j"jjR7&RQ;h2
RRRR8CMRMoCC0sNC(Rz;R

R-RR-VRQR85N8ss_CRo2sHCo#s0CR7q7)#RkHRMoB
piRRRRzR4.RH:RVNR58_8ss2CoRMoCC0sNCR
RRRRRRsRbF#OC#BR5pRi,q)772CRLo
HMRRRRRRRRRRRRH5VRBRpi=4R''MRN8pRBiP'CC2M0RC0EMR
RRRRRRRRRRRRRR8RN_osCRR<=q)7758N8s8IH04E-RI8FMR0Fj
2;RRRRRRRRRRRRCRM8H
V;RRRRRRRRCRM8bOsFC;##
RRRR8CMRMoCC0sNC4Rz.
;
RRRRzR4d:VRHRF5M08RN8ss_CRo2oCCMsCN0
RRRRRRRRRRRR_N8sRCo<q=R757)Ns88I0H8ER-48MFI0jFR2R;
RCRRMo8RCsMCNR0Cz;4d
R
RR.Rzn:RRRRHV5k8F0C_soo2RCsMCN
0CRRRRRRRRbOsFCR##5pmBiF,Rks0_CRo2LHCoMR
RRRRRRRRRRVRHRB5mp=iRR''4R8NMRpmBiP'CC2M0RC0EMR
RRRRRRRRRRRRRRmR7z<aR=kRF0C_soH5I8-0E4FR8IFM0R;j2
RRRRRRRRRRRR8CMR;HV
RRRRRRRR8CMRFbsO#C#;R
RRMRC8CRoMNCs0zCR.
n;
RRRRR--tCCMsCN0RC0ERD#CCRO0DHFoOR
RR4RzcRR:VRFsHMRHRlMk_DOCD8#_CRCb8MFI0jFRRMoCC0sNCR
RR-R-RHAkDF8Rkk0b0MRCNCLDRD#CCRO0DHFoOR
RRRRRR-R-RRQV58N8s8IH0>ERR246RM8F'k0R#1CRpRQBODCD#R
RRRRRR Rm4:nRRRHV58N8s8IH0>ERR246RMoCC0sNCR
RRRRRRRRRRRRRRkRF0M_C5RH2<'=R4I'RERCM5_N8s5CoNs88I0H8ER-48MFI06FR2RR=HC2RDR#C';j'
RRRRRRRR8CMRMoCC0sNC Rm4
n;RRRRRRRR-Q-RVNR58I8sHE80R6>R2hRq7NR58I8sHE80RR<=4R62kR#C1BpQRDOCDR#
RRRRRmRR R46:VRHR85N8HsI8R0E=6R42CRoMNCs0RC
RRRRRRRRRRRRR0RRlNb_858sHg25RI8FMR0Fj<2R=mRhaF5OM#P_0D8_FOoH_OPC05FsH4,RjR22XRm)Ns8_CNo58I8sHE80-84RF0IMF2R6;R
RRRRRRRRRRRRRRqR1h47_6RR:17qh4bjRFRs0lRNb5=qR>lR0b8_N8Hs5225j,RRA=0>RlNb_858sH4252B,RRR=>0_lbNs8855H2.R2,7>R=Rb0l_8N8s25H5,d2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR >R=Rb0l_8N8s25H5,c2R=wR>lR0b8_N8Hs52256,RRt=0>RlNb_858sHn252],RRR=>0_lbNs8855H2(R2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRQ>R=Rb0l_8N8s25H5,U2R=KR>lR0b8_N8Hs5225g,RRZ=F>RkC0_M25H2R;
RRRRRCRRMo8RCsMCNR0Cm6 4;R
RRRRRR Rm4:cRRRHV58N8s8IH0=ERR24cRMoCC0sNCR
RRRRRRRRRRRRRRlR0b8_N8Hs52R5U8MFI0jFR2=R<Rahm5MOFP0_#8F_Do_HOP0COFHs5,2Rg2mRX)8RN_osC58N8s8IH04E-RI8FMR0F6
2;RRRRRRRRRRRRRRRR17qh_R4c:qR1hj74RsbF0NRlbqR5RR=>0_lbNs8855H2jR2,A>R=Rb0l_8N8s25H5,42R=BR>lR0b8_N8Hs5225.,RR7=0>RlNb_858sHd252R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR =0>RlNb_858sHc252w,RRR=>0_lbNs8855H26R2,t>R=Rb0l_8N8s25H5,n2R=]R>lR0b8_N8Hs5225(,RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRQ=0>RlNb_858sHU252K,RRR=>',4'R=ZR>kRF0M_C52H2;R
RRRRRRMRC8CRoMNCs0mCR ;4c
RRRRRRRR4m dRR:H5VRNs88I0H8ERR=4Rd2oCCMsCN0
RRRRRRRRRRRRRRRRb0l_8N8s25H58(RF0IMF2RjRR<=h5maOPFM_8#0_oDFHPO_CFO0s,5HR2U2R)XmR_N8s5CoNs88I0H8ER-48MFI06FR2R;
RRRRRRRRRRRRR1RRq_h74:dRRh1q7RURb0FsRblNRR5q=0>RlNb_858sHj252A,RRR=>0_lbNs8855H24R2,B>R=Rb0l_8N8s25H5,.2R=7R>lR0b8_N8Hs5225d,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR= R>lR0b8_N8Hs5225c,RRw=0>RlNb_858sH6252t,RRR=>0_lbNs8855H2nR2,]>R=Rb0l_8N8s25H5,(2RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR=ZR>kRF0M_C52H2;R
RRRRRRMRC8CRoMNCs0mCR ;4d
RRRRRRRR4m .RR:H5VRNs88I0H8ERR=4R.2oCCMsCN0
RRRRRRRRRRRRRRRRb0l_8N8s25H58nRF0IMF2RjRR<=h5maOPFM_8#0_oDFHPO_CFO0s,5HR2(2R)XmR_N8s5CoNs88I0H8ER-48MFI06FR2R;
RRRRRRRRRRRRR1RRq_h74:.RRh1q7RURb0FsRblNRR5q=0>RlNb_858sHj252A,RRR=>0_lbNs8855H24R2,B>R=Rb0l_8N8s25H5,.2R=7R>lR0b8_N8Hs5225d,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR= R>lR0b8_N8Hs5225c,RRw=0>RlNb_858sH6252t,RRR=>0_lbNs8855H2nR2,]>R=R''4,RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRZ=F>RkC0_M25H2R;
RRRRRCRRMo8RCsMCNR0Cm. 4;R
RRRRRR Rm4:4RRRHV58N8s8IH0=ERR244RMoCC0sNCR
RRRRRRRRRRRRRRlR0b8_N8Hs52R568MFI0jFR2=R<Rahm5MOFP0_#8F_Do_HOP0COFHs5,2Rn2mRX)8RN_osC58N8s8IH04E-RI8FMR0F6
2;RRRRRRRRRRRRRRRR17qh_R44:qR1hR7nRsbF0NRlbqR5RR=>0_lbNs8855H2jR2,A>R=Rb0l_8N8s25H5,42R=BR>lR0b8_N8Hs5225.,RR7=0>RlNb_858sHd252R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR =0>RlNb_858sHc252w,RRR=>0_lbNs8855H26R2,Z>R=R0Fk_5CMH;22
RRRRRRRR8CMRMoCC0sNC Rm4
4;RRRRRRRRmj 4RH:RVNR58I8sHE80R4=Rjo2RCsMCN
0CRRRRRRRRRRRRRRRR0_lbNs8855H2cFR8IFM0RRj2<h=RmOa5F_MP#_08DHFoOC_POs0F5RH,6R22XRm)Ns8_CNo58I8sHE80-84RF0IMF2R6;R
RRRRRRRRRRRRRRqR1h47_jRR:17qhnbRRFRs0lRNb5=qR>lR0b8_N8Hs5225j,RRA=0>RlNb_858sH4252B,RRR=>0_lbNs8855H2.R2,7>R=Rb0l_8N8s25H5,d2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR >R=Rb0l_8N8s25H5,c2R=wR>4R''Z,RRR=>F_k0CHM52
2;RRRRRRRRCRM8oCCMsCN0R4m jR;
RRRRRmRR RgR:VRHR85N8HsI8R0E=2RgRMoCC0sNCR
RRRRRRRRRRRRRRlR0b8_N8Hs52R5d8MFI0jFR2=R<Rahm5MOFP0_#8F_Do_HOP0COFHs5,2Rc2mRX)8RN_osC58N8s8IH04E-RI8FMR0F6
2;RRRRRRRRRRRRRRRR17qh_:gRRh1q7RcRRsbF0NRlbqR5RR=>0_lbNs8855H2jR2,A>R=Rb0l_8N8s25H5,42R=BR>lR0b8_N8Hs5225.,RR7=0>RlNb_858sHd252R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRZ=F>RkC0_M25H2R;
RRRRRCRRMo8RCsMCNR0Cm; g
RRRRRRRRUm RRR:H5VRNs88I0H8ERR=Uo2RCsMCN
0CRRRRRRRRRRRRRRRR0_lbNs8855H2.FR8IFM0RRj2<h=RmOa5F_MP#_08DHFoOC_POs0F5RH,dR22XRm)Ns8_CNo58I8sHE80-84RF0IMF2R6;R
RRRRRRRRRRRRRRqR1hU7_R1:Rqch7RbRRFRs0lRNb5=qR>lR0b8_N8Hs5225j,RRA=0>RlNb_858sH4252B,RRR=>0_lbNs8855H2.R2,7>R=R''4,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR=ZR>kRF0M_C52H2;R
RRRRRRMRC8CRoMNCs0mCR 
U;RRRRRRRRmR (RH:RVNR58I8sHE80R(=R2CRoMNCs0RC
RRRRRRRRRRRRR0RRlNb_858sH425RI8FMR0Fj<2R=mRhaF5OM#P_0D8_FOoH_OPC05FsH.,R2X2RmN)R8C_so85N8HsI8-0E4FR8IFM0R;62
RRRRRRRRRRRRRRRRh1q7R_(:qR1hR7.RFRbsl0RN5bRq>R=Rb0l_8N8s25H5,j2R=AR>lR0b8_N8Hs52254,RRZ=F>RkC0_M25H2R;
RRRRRCRRMo8RCsMCNR0Cm; (
RRRRRRRRnm RRR:H5VRNs88I0H8ERR=no2RCsMCN
0CRRRRRRRRRRRRRRRRF_k0CHM52=R<R''4RCIEMNR58C_so256RO=RF_MP#_08DHFoOC_POs0F54H,225j2DRC#'CRj
';RRRRRRRRCRM8oCCMsCN0Rnm ;R
RR-R-RRQV58N8s8IH0<ER=2R6RRMFFbk0kC0RMDNLCCR#D0CORoDFHMORCCC88RR/lRNb8CHsO$0DRR0F)'qv#8RN8#sC#HRDM
C#RRRRRRRRmR 6:VRHR85N8HsI8R0E<6=R2CRoMNCs0RC
RRRRRRRRRRRRRFRRkC0_M25HRR<=';4'
RRRRRRRR8CMRMoCC0sNC Rm6
;
RRRR-Q-RVNR58I8sHE80Rg>R2#RkCuRW 0jRFCR8OCF8R8N8s#C#R0LH#RRn0FEskRoEgMRN8uRW 04RFCR8OCF8R0LH#jR4RR+
RRRRRWRR R4j:VRHR85N8HsI8R0E>2RgRMoCC0sNCR
RRRRRRRRRRRRRRbRICCj_M25HRR<='R4'IMECR85N_osC58URF0IMF2R6RO=RF_MP#_08DHFoOC_POs0F5.H,jd25RI8FMR0FjR22CCD#R''j;R
RRRRRRRRRRRRRRbRICC4_M25HRR<='R4'IMECR85N_osC58N8s8IH04E-RI8FMR0Fg=2RRMOFP0_#8F_Do_HOP0COFHs5,2.j58N8s8IH0nE-RI8FMR0FcR22CCD#R''j;R
RRRRRRRRRRMRC8CRoMNCs0WCR ;4j
RRRRR--Q5VRNs88I0H8ERR=UsRFRRg2kR#CWju RR0F8FCO8NCR8C8s#L#RHR0#nER0soFkE
RgRRRRRRRRWR gRH:RV5R5Ns88I0H8ERR=Um2R)NR58I8sHE80Rg=R2o2RCsMCN
0CRRRRRRRRRRRRRRRRIjbC_5CMH<2R=4R''ERIC5MRNs8_CNo58I8sHE80-84RF0IMF2R6RH=R2DRC#'CRj
';RRRRRRRRRRRRRRRRI4bC_5CMH<2R=4R''R;
RRRRRRRRRCRRMo8RCsMCNR0CW; g
RRRRR--Q5VRNs88I0H8ERR=(k2R#WCRuR j08FRC8OFCER0C0RnE8RN8#sC#HRL0RR&W4u RR0F8FCO80CRE(CR0NER8C8s#L#RHR0
RRRRRWRR R(R:VRHR85N8HsI8R0E=2R(RMoCC0sNCR
RRRRRRRRRRRRRRbRICCj_M25HRR<='R4'IMECR85N_osC5R62=FROM#P_0D8_FOoH_OPC05FsH2,.52j2R#CDCjR''R;
RRRRRRRRRRRRRIRRb_C4CHM52=R<R''4RCIEMNR58C_so25nRO=RF_MP#_08DHFoOC_POs0F5.H,22542DRC#'CRj
';RRRRRRRRCRM8oCCMsCN0R(W ;R
RR-R-RRQV58N8s8IH0=ERRRn2kR#CWju RR0F8FCO80CREnCR0NER8C8s#L#RHR0
RRRRRWRR RnR:VRHR85N8HsI8R0E=2RnRMoCC0sNCR
RRRRRRRRRRRRRRbRICCj_M25HRR<='R4'IMECR85N_osC5R62=FROM#P_0D8_FOoH_OPC05FsH2,452j2R#CDCjR''R;
RRRRRRRRRRRRRIRRb_C4CHM52=R<R''4;R
RRRRRRMRC8CRoMNCs0WCR 
n;RRRR-Q-RVNR58I8sHE80RR<=6M2RFsRIHR0CCLMND#CRCODC0FRDoRHOM8CCCR8
RRRRRWRR R6R:VRHR85N8HsI8R0E<6=R2CRoMNCs0RC
RRRRRRRRRRRRRIRRb_CjCHM52=R<R''4;R
RRRRRRRRRRRRRRbRICC4_M25HRR<=';4'
RRRRRRRR8CMRMoCC0sNC RW6
;
RRRRCRM8oCCMsCN0Rcz4;R

RzRR.:6RRRHV50MFRk8F0C_soo2RCsMCN
0CRRRRRRRRz44(:sRbF#OC#FR5ks0_C
o2RRRRRRRRLHCoMR
RRRRRRRRRRmR7z<aR=kRF0C_soH5I8-0E4FR8IFM0R;j2
RRRRRRRR8CMRFbsO#C#R(z44R;
RCRRMo8RCsMCNR0Cz;.6
R
RR-R-RMtCC0sNCER0CqR)vCRODRD#IEH0RH0s-N#00
C#RRRRzR46:FRVsRRHHMMRkOl_C#DD_C8CbFR8IFM0RojRCsMCN
0CRRRRRRRRzR4(:FRVsRR[HMMRkOl_C#DD_8IHCFR8IFM0RojRCsMCN
0CRRRRRRRRRRRRzv)q:BR) Xd.cRR
RRRRRRRRRRRRRbRRFRs0lRNb5j7QRR=>HsM_C5o5[2*c27,RQ=4R>MRH_osC5*5[c42+27,RQ=.R>MRH_osC5*5[c.2+27,RQ=dR>MRH_osC5*5[cd2+2t,R1=)R>4R''
,RRRRRRRRRRRRRRRRRRRRRRRRRR7Rqj>R=RIDF_8N8s25j,7Rq4>R=RIDF_8N8s254,7Rq.>R=RIDF_8N8s25.,7Rqd>R=RIDF_8N8s25d,7Rqc>R=RIDF_8N8s25c,-R
-RRRRRRRRRRRRRRRRRRRRRRRRWRR)R h=W>R W,RuR j=I>Rb_CjCHM52W,RuR 4=I>Rb_C4CHM52B,Ri>R=RahmRiBp,RR
RRRRRRRRRRRRRRRRRRRRRRRRR W)h>R=R,W R Wuj>R=RCIbjM_C5,H2R Wu4>R=RCIb4M_C5,H2RRBi=B>RpRi,
RRRRRRRRRRRRRRRRRRRRRRRR7RRm=jR>kRF0k_L#,5H5c[*2R2,7Rm4=F>RkL0_kH#5,*5[c42+27,Rm=.R>kRF0k_L#,5H5c[*22+.,mR7d>R=R0Fk_#Lk55H,[2*c+2d2;R
RRRRRRRRRRRRRRkRF0C_so[55*2c2RR<=F_k0L5k#H[,5*2c2RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_so[55*+c24<2R=kRF0k_L#,5H5c[*22+4RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_so[55*+c2.<2R=kRF0k_L#,5H5c[*22+.RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_so[55*+c2d<2R=kRF0k_L#,5H5c[*22+dRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRMRC8CRoMNCs0zCR4
(;RRRRRRRRCRM8oCCMsCN0R6z4;-

-zRR.:URRRHV5k8F0C_soo2RCsMCN
0C-R-RRRRRR4RznRR:VRFsHMRHRlMk_DOCD8#_CRCb8MFI0jFRRMoCC0sNC-
-RRRRRRRRzR4U:FRVsRR[HMMRkOl_C#DD_8IHCFR8IFM0RojRCsMCN
0C-R-RRRRRRRRRR)RzqRv:)dB .RXc
R--RRRRRRRRRRRRRbRRFRs0lRNb5j7QRR=>HsM_C5o5[2*c27,RQ=4R>MRH_osC5*5[c42+27,RQ=.R>MRH_osC5*5[c.2+27,RQ=dR>MRH_osC5*5[cd2+2-,
-RRRRRRRRRRRRRRRRRRRRRRRRqRR7=jR>FRDI8_N8js52q,R7=4R>FRDI8_N84s52q,R7=.R>FRDI8_N8.s52q,R7=dR>FRDI8_N8ds52q,R7=cR>FRDI8_N8cs52-,
-RRRRRRRRRRRRRRRRRRRRRRRRWRR)R h=W>R W,RuR j=I>Rb_CjCHM52W,RuR 4=I>Rb_C4CHM52B,Ri>R=RahmRiBp,-R
-RRRRRRRRRRRRRRRRRRRRRRRRTRR7Rmj=F>RkL0_kH#5,*5[c,22RmT74>R=R0Fk_#Lk55H,[2*c+,42RmT7.>R=R0Fk_#Lk55H,[2*c+,.2RmT7d>R=R0Fk_#Lk55H,[2*c+2d2;-
-RRRRRRRRRRRRRRRRF_k0s5Co5c[*2<2R=kRF0k_L#,5H5c[*2I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';-R-RRRRRRRRRRRRRRkRF0C_so[55*+c24<2R=kRF0k_L#,5H5c[*22+4RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;-
-RRRRRRRRRRRRRRRRF_k0s5Co5c[*22+.RR<=F_k0L5k#H[,5*+c2.I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';-R-RRRRRRRRRRRRRRkRF0C_so[55*+c2d<2R=kRF0k_L#,5H5c[*22+dRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;-
-RRRRRRRRRRRRCRM8oCCMsCN0RUz4;-
-RRRRRCRRMo8RCsMCNR0Cz;4n
R--RCRRMo8RCsMCNR0Cz;.U
-
-RRRRRURkRH:RV8R5F_k0s2CoRMoCC0sNC-
-RRRRRRRRRmR7z<aR=kRF0C_soH5I8-0E4FR8IFM0R;j2
R--R8CMRMoCC0sNCURk;R
RRRRRRRRRRRRRR
RRCRM8NEsOHO0C0CksRONsE
j;
