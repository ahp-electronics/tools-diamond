-- ---------------------------------------------------------------------------
--
-- Name : ER1.vhd
--
-- Description:
--
--    This module is where the ER1 register implemented. ER1 and ER2 registers
--    can be registers implemented in Lattice FPGAs using normal FPGA's
--    programmable logic resources.  Once they are implemented, they can be
--    accessed as if they are JTAG data registers through the FPGA JTAG port.
--    In order to accessing these registers, JTAG instructions ER1(0x32) or
--    ER2(0x38) needs to be written to the JTAG IR register for enabling the
--    ER1/ER2 accessing logic.  The ER1 or ER2 accessing logic can only be
--    enabled one at a time.  Once they are enabled, they will be disabled if
--    another JTAG instruction is written into the JTAG instruction register.
--    The registers allow dynamically accessing the FPGA internal information
--    even when the device is running.  Therefore, they are very useful for some
--    of the IP cores.  In order to let ER1/ER2 registers shared by multiple IP
--    cores or other designs, there is a ER1/ER2 structure patterned by Lattice.
--    The ER1/ER2 structure allows only one ER1 register but more than one ER2
--    registers in an FPGA device.  Please refer to the related document for
--    this patterned ER1/ER2 structure.
--
-- $Log: er1.vhd,v $
-- Revision 1.3  2005-03-17 17:19:36-08  jhsin
-- Added ER1, ER2 attributes to turn on the ER1, ER2 fuses in XP.
--
-- Revision 1.2  2004-10-08 16:17:50-07  jhsin
-- Added port "ISPTRACY_ER2_TDO" for reading back ispTRACY er2 registers.
--
-- Revision 1.1  2004-09-09 11:41:12-07  jhsin
-- Moved JTAGB instantiation from the top level module (spitop.vhd)
-- to ER1 module.  Now the ER1 module is a common module and can
-- be used for SPI Serial FLASH Programmer, ispTRACY and other IPs.
--
-- Revision 1.0  2004-08-03 18:35:56-07  jhsin
-- Initial revision
--
--
-- $Header: \\\\hqfs2\\ip\040cores\\rcs\\hqfs2\\ip\040cores\\rcswork\\isptracy\\VHDL\\Implementation\\er1.vhd,v 1.3 2005-03-17 17:19:36-08 jhsin Exp $
--
-- Copyright (C) 2004 Lattice Semiconductor Corp.  All rights reserved.
--
-- ---------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

entity ER1 is
   port (
      JTCK             : out std_logic;
      JTDI             : out std_logic;
      JSHIFT           : out std_logic;
      JUPDATE          : out std_logic;
      JRSTN            : out std_logic;
      JCE2             : out std_logic;
      JRTI2            : out std_logic;
      ER2_TDO          : in  std_logic_vector(14 downto 0);
      ISPTRACY_ER2_TDO : in  std_logic;
      IP_ENABLE        : out std_logic_vector(14 downto 0);
      ISPTRACY_ENABLE  : out std_logic;
      CONTROL_DATAN    : out std_logic
   );
end ER1;

architecture ER1_a of ER1 is

   component JTAGB
      port (
         JTCK    : out std_logic;
         JRTI1   : out std_logic;
         JRTI2   : out std_logic;
         JTDI    : out std_logic;
         JSHIFT  : out std_logic;
         JUPDATE : out std_logic;
         JRSTN   : out std_logic;
         JCE1    : out std_logic;
         JCE2    : out std_logic;
         JTDO1   : in  std_logic;
         JTDO2   : in  std_logic
      );
   end component;

   component TYPEA
      port (
         CLK        : in  std_logic;
         RESET_N    : in  std_logic;
         CLKEN      : in  std_logic;
         TDI        : in  std_logic;
         TDO        : out std_logic;
         DATA_OUT   : out std_logic;
         DATA_IN    : in  std_logic;
         CAPTURE_DR : in  std_logic;
         UPDATE_DR  : in  std_logic
      );
   end component;

   component TYPEB
      port (
         CLK        : in  std_logic;
         RESET_N    : in  std_logic;
         CLKEN      : in  std_logic;
         TDI        : in  std_logic;
         TDO        : out std_logic;
         DATA_IN    : in  std_logic;
         CAPTURE_DR : in  std_logic
      );
   end component;

   signal tck       : std_logic;
   signal tdi       : std_logic;
   signal shiftDr   : std_logic;
   signal updateDr  : std_logic;
   signal resetN    : std_logic;
   signal enableEr1 : std_logic;
   signal tdoEr1    : std_logic;
   signal tdoEr2    : std_logic;

   signal controlDataNBit     : std_logic;
   signal ispTracyEnableBit   : std_logic;
   signal encodedIpEnableBits : std_logic_vector(3 downto 0);
   signal er1TdiBit           : std_logic_vector(9 downto 0);
   signal captureDrER1        : std_logic;

   attribute ER1 : string; 
   attribute ER1 of DEDICATE_LOGIC : label is "ENABLED";
   attribute ER2 : string; 
   attribute ER2 of DEDICATE_LOGIC : label is "ENABLED";

begin

   JTCK    <= tck;
   JTDI    <= tdi;
   JSHIFT  <= shiftDr;
   JUPDATE <= updateDr;
   JRSTN   <= resetN;

   DEDICATE_LOGIC : JTAGB
   port map (
      JTCK    => tck,
      JRTI1   => open,
      JRTI2   => JRTI2,
      JTDI    => tdi,
      JSHIFT  => shiftDr,
      JUPDATE => updateDr,
      JRSTN   => resetN,
      JCE1    => enableEr1,
      JCE2    => JCE2,
      JTDO1   => tdoEr1,
      JTDO2   => tdoEr2
   );

   tdoEr1 <= er1TdiBit(0);

   BIT0 : TYPEB
   port map (
      CLK        => tck,
      RESET_N    => resetN,
      CLKEN      => enableEr1,
      TDI        => er1TdiBit(1),
      TDO        => er1TdiBit(0),
      DATA_IN    => '0',
      CAPTURE_DR => captureDrER1
   );

   BIT1 : TYPEB
   port map (
      CLK        => tck,
      RESET_N    => resetN,
      CLKEN      => enableEr1,
      TDI        => er1TdiBit(2),
      TDO        => er1TdiBit(1),
      DATA_IN    => '0',
      CAPTURE_DR => captureDrER1
   );

   BIT2 : TYPEB
   port map (
      CLK        => tck,
      RESET_N    => resetN,
      CLKEN      => enableEr1,
      TDI        => er1TdiBit(3),
      TDO        => er1TdiBit(2),
      DATA_IN    => '1',
      CAPTURE_DR => captureDrER1
   );

   BIT3 : component TYPEA
   port map (
      CLK        => tck,
      RESET_N    => resetN,
      CLKEN      => enableEr1,
      TDI        => er1TdiBit(4),
      TDO        => er1TdiBit(3),
      DATA_OUT   => controlDataNBit,
      DATA_IN    => controlDataNBit,
      CAPTURE_DR => captureDrER1,
      UPDATE_DR  => updateDr
   );

   CONTROL_DATAN <= controlDataNBit;

   BIT4 : component TYPEA
   port map (
      CLK        => tck,
      RESET_N    => resetN,
      CLKEN      => enableEr1,
      TDI        => er1TdiBit(5),
      TDO        => er1TdiBit(4),
      DATA_OUT   => ispTracyEnableBit,
      DATA_IN    => ispTracyEnableBit,
      CAPTURE_DR => captureDrER1,
      UPDATE_DR  => updateDr
   );

   ISPTRACY_ENABLE <= ispTracyEnableBit;

   BIT5_BIT8 : for bit_index in 5 to 8 generate
   begin
      BIT_N : component TYPEA
      port map (
         CLK        => tck,
         RESET_N    => resetN,
         CLKEN      => enableEr1,
         TDI        => er1TdiBit(bit_index + 1),
         TDO        => er1TdiBit(bit_index),
         DATA_OUT   => encodedIpEnableBits(bit_index - 5),
         DATA_IN    => encodedIpEnableBits(bit_index - 5),
         CAPTURE_DR => captureDrER1,
         UPDATE_DR  => updateDr
      );
   end generate BIT5_BIT8;

   er1TdiBit(9) <= tdi;

   captureDrER1  <= not shiftDr and enableEr1;

   DECODE : process (encodedIpEnableBits, ER2_TDO) is
   begin
      case encodedIpEnableBits is
         when "0000" =>
            IP_ENABLE <= "000000000000000";
            tdoEr2    <= ISPTRACY_ER2_TDO;
         when "0001" =>
            IP_ENABLE <= "000000000000001";
            tdoEr2    <= ER2_TDO(0);
         when "0010" =>
            IP_ENABLE <= "000000000000010";
            tdoEr2    <= ER2_TDO(1);
         when "0011" =>
            IP_ENABLE <= "000000000000100";
            tdoEr2    <= ER2_TDO(2);
         when "0100" =>
            IP_ENABLE <= "000000000001000";
            tdoEr2    <= ER2_TDO(3);
         when "0101" =>
            IP_ENABLE <= "000000000010000";
            tdoEr2    <= ER2_TDO(4);
         when "0110" =>
            IP_ENABLE <= "000000000100000";
            tdoEr2    <= ER2_TDO(5);
         when "0111" =>
            IP_ENABLE <= "000000001000000";
            tdoEr2    <= ER2_TDO(6);
         when "1000" =>
            IP_ENABLE <= "000000010000000";
            tdoEr2    <= ER2_TDO(7);
         when "1001" =>
            IP_ENABLE <= "000000100000000";
            tdoEr2    <= ER2_TDO(8);
         when "1010" =>
            IP_ENABLE <= "000001000000000";
            tdoEr2    <= ER2_TDO(9);
         when "1011" =>
            IP_ENABLE <= "000010000000000";
            tdoEr2    <= ER2_TDO(10);
         when "1100" =>
            IP_ENABLE <= "000100000000000";
            tdoEr2    <= ER2_TDO(11);
         when "1101" =>
            IP_ENABLE <= "001000000000000";
            tdoEr2    <= ER2_TDO(12);
         when "1110" =>
            IP_ENABLE <= "010000000000000";
            tdoEr2    <= ER2_TDO(13);
         when "1111" =>
            IP_ENABLE <= "100000000000000";
            tdoEr2    <= ER2_TDO(14);
         when others =>
            IP_ENABLE <= "000000000000000";
            tdoEr2    <= '0';
      end case;
   end process DECODE;

end ER1_a;
-- ---------------------------------------------------------------------------
--
-- Name : SPIPROG.vhd
--
-- Description:
--
--    This module contains the ER2 regsiters of SPI Serial FLASH programmer IP
--    core.  There are only three ER2 registers, one control register and two
--    data registers, in this IP core.  The control register is a 8-bit wide
--    register for selecting which data register will be accessed when the
--    Control/Data# bit in ER1 register is low.  Data register 0 is a readonly
--    ID register.  It is composed of three register fields -- an 8-bit
--    "implementer", a 16-bit "IP_functionality", and a 12-bit "revision".
--    Data register 1 is a variable length register for sending commands to or
--    receiving readback data from the SPI Serial FLASH device.
--
-- $Log: spiprog.vhd,v $
-- Revision 1.3  2004-10-08 16:19:46-07  jhsin
-- Added 1-bit DR2 register for tri-stating outputs after SPI programming completed.
--
-- Revision 1.2  2004-09-09 11:43:26-07  jhsin
-- 1. Reduced the the ID register (DR0) length from 36 bits to 8 bits.
-- 2. Same as TYPEA and TYPEB modules, use falling edge clock
--    for all TCK Flip-Flops.
--
-- Revision 1.1  2004-08-12 13:22:05-07  jhsin
-- Added 7 delay Flip-Flops so that the DR1 readback data from SPI Serial FLASH is in the byte boundary.
--
-- Revision 1.0  2004-08-03 18:35:56-07  jhsin
-- Initial revision
--
--
-- $Header: \\\\hqfs2\\ip\040cores\\rcs\\hqfs2\\ip\040cores\\rcswork\\isptracy\\VHDL\\Implementation\\spiprog.vhd,v 1.3 2004-10-08 16:19:46-07 jhsin Exp $
--
-- Copyright (C) 2004 Lattice Semiconductor Corp.  All rights reserved.
--
-- ---------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

entity SPIPROG is
   port (
      JTCK           : in  std_logic;
      JTDI           : in  std_logic;
      JTDO2          : out std_logic;
      JSHIFT         : in  std_logic;
      JUPDATE        : in  std_logic;
      JRSTN          : in  std_logic;
      JCE2           : in  std_logic;
      SPIPROG_ENABLE : in  std_logic;
      CONTROL_DATAN  : in  std_logic;
      SPI_C          : out std_logic;
      SPI_D          : out std_logic;
      SPI_SN         : out std_logic;
      SPI_Q          : in  std_logic
   );
end SPIPROG;

architecture SPIPROG_a of SPIPROG is

   component TYPEA
      port (
         CLK        : in  std_logic;
         RESET_N    : in  std_logic;
         CLKEN      : in  std_logic;
         TDI        : in  std_logic;
         TDO        : out std_logic;
         DATA_OUT   : out std_logic;
         DATA_IN    : in  std_logic;
         CAPTURE_DR : in  std_logic;
         UPDATE_DR  : in  std_logic
      );
   end component;

   component TYPEB
      port (
         CLK        : in  std_logic;
         RESET_N    : in  std_logic;
         CLKEN      : in  std_logic;
         TDI        : in  std_logic;
         TDO        : out std_logic;
         DATA_IN    : in  std_logic;
         CAPTURE_DR : in  std_logic
      );
   end component;

   signal er2Cr_enable  : std_logic;
   signal er2Dr0_enable : std_logic;
   signal er2Dr1_enable : std_logic;
   signal er2Dr2_enable : std_logic;

   signal tdo_er2Cr  : std_logic;
   signal tdo_er2Dr0 : std_logic;
   signal tdo_er2Dr1 : std_logic;
   signal tdo_er2Dr2 : std_logic;

   signal encodedDrSelBits : std_logic_vector(7 downto 0);
   signal er2CrTdiBit      : std_logic_vector(8 downto 0);
   signal er2Dr0TdiBit     : std_logic_vector(8 downto 0);

   signal captureDrER2 : std_logic;
   signal spi_s        : std_logic;
   signal spi_q_dly    : std_logic_vector(6 downto 0);

   signal spi_c_i  : std_logic;
   signal spi_d_i  : std_logic;
   signal spi_sn_i : std_logic;

   signal triStateOutput : std_logic;

   signal ip_functionality_id : std_logic_vector(7 downto 0);

begin

   ------ Control Register 0 ------

   er2Cr_enable <= JCE2 and SPIPROG_ENABLE and CONTROL_DATAN;

   tdo_er2Cr <= er2CrTdiBit(0);

   CR_BIT0_BIT7 : for bit_index in 0 to 7 generate
   begin
      BIT_N : component TYPEA
      port map (
         CLK        => JTCK,
         RESET_N    => JRSTN,
         CLKEN      => er2Cr_enable,
         TDI        => er2CrTdiBit(bit_index + 1),
         TDO        => er2CrTdiBit(bit_index),
         DATA_OUT   => encodedDrSelBits(bit_index),
         DATA_IN    => encodedDrSelBits(bit_index),
         CAPTURE_DR => captureDrER2,
         UPDATE_DR  => JUPDATE
      );
   end generate CR_BIT0_BIT7;

   er2CrTdiBit(8) <= JTDI;

   ------ Data Register 0 ------

   er2Dr0_enable <= '1' when (JCE2 = '1') and (SPIPROG_ENABLE = '1') and (CONTROL_DATAN = '0') and (encodedDrSelBits = "00000000") else
                    '0';

   tdo_er2Dr0 <= er2Dr0TdiBit(0);

   ip_functionality_id <= "00000001";  -- SPI Serial FLASH Programmer (0x01)

   DR0_BIT0_BIT7 : for bit_index in 0 to 7 generate
   begin
      BIT_N : TYPEB
      port map (
         CLK        => JTCK,
         RESET_N    => JRSTN,
         CLKEN      => er2Dr0_enable,
         TDI        => er2Dr0TdiBit(bit_index + 1),
         TDO        => er2Dr0TdiBit(bit_index),
         DATA_IN    => ip_functionality_id(bit_index),
         CAPTURE_DR => captureDrER2
      );
   end generate DR0_BIT0_BIT7;

   er2Dr0TdiBit(8) <= JTDI;

   ------ Data Register 1 ------

   er2Dr1_enable <= '1' when (JCE2 = '1') and (JSHIFT = '1') and (SPIPROG_ENABLE = '1') and (CONTROL_DATAN = '0') and (encodedDrSelBits = "00000001") else
                    '0';

   spi_c_i <= not (JTCK and er2Dr1_enable and spi_s);

   spi_d_i <= JTDI and er2Dr1_enable;

   SPI_S_Proc : process (JTCK, JRSTN)
   begin
      if (JRSTN='0') then
         spi_s <= '0';
      elsif falling_edge(JTCK) then
         if (JUPDATE = '1') then
            spi_s <= '0';
         else
            spi_s <= er2Dr1_enable;
         end if;
      end if;
   end process SPI_S_Proc;

   spi_sn_i <= not spi_s;

   SPI_Q_Proc : process (JTCK, JRSTN)
   begin
      if (JRSTN='0') then
         spi_q_dly <= (others => '0');
      elsif falling_edge(JTCK) then
         if (er2Dr1_enable = '1') then
            spi_q_dly  <= spi_q_dly(5 downto 0) & SPI_Q;
         end if;
      end if;
   end process SPI_Q_Proc;

   tdo_er2Dr1 <= spi_q_dly(6);

   ------ Data Register 2 ------

   er2Dr2_enable <= '1' when (JCE2 = '1') and (SPIPROG_ENABLE = '1') and (CONTROL_DATAN = '0') and (encodedDrSelBits = "00000010") else
                    '0';

   DR2_BIT0 : TYPEA
      port map (
         CLK        => JTCK,
         RESET_N    => JRSTN,
         CLKEN      => er2Dr2_enable,
         TDI        => JTDI,
         TDO        => tdo_er2Dr2,
         DATA_OUT   => triStateOutput,
         DATA_IN    => triStateOutput,
         CAPTURE_DR => captureDrER2,
         UPDATE_DR  => JUPDATE
      );

   ------ OUTPUT TRI-STATE CONTROL ------

   SPI_C  <=  spi_c_i when (triStateOutput = '0') else 'Z';
   SPI_D  <=  spi_d_i when (triStateOutput = '0') else 'Z';
   SPI_SN <= spi_sn_i when (triStateOutput = '0') else 'Z';

   ------ JTDO2 MUX ------

   JTDO2 <= tdo_er2Cr when (CONTROL_DATAN = '1') else
            tdo_er2Dr0 when (CONTROL_DATAN = '0') and (encodedDrSelBits = "00000000") else
            tdo_er2Dr1 when (CONTROL_DATAN = '0') and (encodedDrSelBits = "00000001") else
            tdo_er2Dr2 when (CONTROL_DATAN = '0') and (encodedDrSelBits = "00000010") else
            '0';

   captureDrER2  <= not JSHIFT and JCE2;

end SPIPROG_a;
-- ---------------------------------------------------------------------------
--
-- Name : TYPEA.vhd
--
-- Description:
--
--    This is one of the two types of cells that are used to create ER1/ER2
--    register bits.
--
-- $Log: typea.vhd,v $
-- Revision 1.3  2004-09-02 15:31:19-07  jhsin
-- Changed all the ispTRACY internal type-A and type-B registers from rising edge
-- registers to falling edge registers.  The write enable and write address signals
-- in the MAPW module are changed as well.  Now the event comparison RAM
-- and trigger RAM are written at the falling edge of TCK.
--
-- Revision 1.2  2002-11-13 18:33:59-08  jhsin
-- The SHIFT_DR_CAPTURE_DR and ENABLE_ER1/2 signals of the
-- dedicate logic JTAG_PORT didn't act as what their names implied.
-- The SHIFT_DR_CAPTURE_DR actually acts as SHIFT_DR.
-- The ENABLE_ER1/2 actually acts as SHIFT_DR_CAPTURE_DR.
-- These had caused a lot of headaches for a long time and now they are
-- fixed by:
-- (1) Use SHIFT_DR_CAPTURE_DR and ENABLE_ER1/2 to create
--     CAPTURE_DR for all typeA, typeB bits in the ER1, ER2 registers.
-- (2) Use ENABLE_ER1 or the enESR, enCSR, enBAR (these 3 signals
--     have the same waveform of ENABLE_ER2) directly to be the CLKEN
--     of all typeA, typeB bits in the ER1, ER2 registers.
-- (3) Modify typea.vhd to use only UPDATE_DR signal for the clock enable
--     of the holding flip-flop.
-- These changes caused ispTracy.vhd and cge.dat changes and the new
-- CGE.exe version will be 1.3.5.
--
-- Revision 1.1  2002-05-01 18:13:51-07  jhsin
-- Added RCS version control header to file. No code changes.
--
-- $Header: \\\\hqfs2\\ip\040cores\\rcs\\hqfs2\\ip\040cores\\rcswork\\isptracy\\VHDL\\Implementation\\typea.vhd,v 1.3 2004-09-02 15:31:19-07 jhsin Exp $
--
-- Copyright (C) 2002 Lattice Semiconductor Corp.  All rights reserved.
--
-- ---------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

entity TYPEA is
   port (
      CLK        : in  std_logic;
      RESET_N    : in  std_logic;
      CLKEN      : in  std_logic;
      TDI        : in  std_logic;
      TDO        : out std_logic;
      DATA_OUT   : out std_logic;
      DATA_IN    : in  std_logic;
      CAPTURE_DR : in  std_logic;
      UPDATE_DR  : in  std_logic
   );
end TYPEA;

architecture TYPEA_a of TYPEA is

   signal tdoInt : std_logic;

begin

   CAPTURE_Proc : process (CLK, RESET_N)
   begin
      if (RESET_N='0') then
         tdoInt <= '0';
      elsif falling_edge(CLK) then
         if (CLKEN='1') then
            if (CAPTURE_DR='0') then
               tdoInt <= TDI;
            else
               tdoInt <= DATA_IN;
            end if;
         end if;
      end if;
   end process CAPTURE_Proc;

   TDO <= tdoInt;

   UPDATE_Proc : process (CLK, RESET_N)
   begin
      if (RESET_N='0') then
         DATA_OUT <= '0';
      elsif falling_edge(CLK) then
         if (UPDATE_DR='1') then
            DATA_OUT <= tdoInt;
         end if;
      end if;
   end process UPDATE_Proc;

end TYPEA_a;

-- ---------------------------------------------------------------------------
--
-- Name : TYPEB.vhd
--
-- Description:
--
--    This is one of the two types of cells that are used to create ER1/ER2
--    register bits.
--
-- $Log: typeb.vhd,v $
-- Revision 1.3  2004-09-02 15:31:18-07  jhsin
-- Changed all the ispTRACY internal type-A and type-B registers from rising edge
-- registers to falling edge registers.  The write enable and write address signals
-- in the MAPW module are changed as well.  Now the event comparison RAM
-- and trigger RAM are written at the falling edge of TCK.
--
-- Revision 1.2  2002-08-01 16:39:33-07  jhsin
-- Modified typeb module to remove redundant DATA_OUT port.
--
-- Revision 1.1  2002-05-01 18:13:51-07  jhsin
-- Added RCS version control header to file. No code changes.
--
-- $Header: \\\\hqfs2\\ip\040cores\\rcs\\hqfs2\\ip\040cores\\rcswork\\isptracy\\VHDL\\Implementation\\typeb.vhd,v 1.3 2004-09-02 15:31:18-07 jhsin Exp $
--
-- Copyright (C) 2002 Lattice Semiconductor Corp.  All rights reserved.
--
-- ---------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

entity TYPEB is
   port (
      CLK        : in  std_logic;
      RESET_N    : in  std_logic;
      CLKEN      : in  std_logic;
      TDI        : in  std_logic;
      TDO        : out std_logic;
      DATA_IN    : in  std_logic;
      CAPTURE_DR : in  std_logic
   );
end TYPEB;

architecture TYPEB_a of TYPEB is

   signal tdoInt : std_logic;

begin

   CAPTURE_Proc : process (CLK, RESET_N)
   begin
      if (RESET_N='0') then
         tdoInt <= '0';
      elsif falling_edge(CLK) then
         if (CLKEN='1') then
            if (CAPTURE_DR='0') then
               tdoInt <= TDI;
            else
               tdoInt <= DATA_IN;
            end if;
         end if;
      end if;
   end process CAPTURE_Proc;

   TDO <= tdoInt;

end TYPEB_a;

