library verilog;
use verilog.vl_types.all;
entity pp_rx_top is
    port(
        rx_clk          : in     vl_logic;
        ebrd_clk        : in     vl_logic;
        rst_rx_clk_n    : in     vl_logic;
        rst_ebrd_clk_n  : in     vl_logic;
        rxd_i           : in     vl_logic_vector(9 downto 0);
        rxd_o           : out    vl_logic_vector(11 downto 0);
        tobist_data1    : out    vl_logic_vector(9 downto 0);
        ls_sync_status  : out    vl_logic;
        cc_re_o         : out    vl_logic;
        cc_we_o         : out    vl_logic;
        loopback        : in     vl_logic;
        signal_detect   : in     vl_logic;
        enable_cgalign  : in     vl_logic;
        udf_comma_a     : in     vl_logic_vector(9 downto 0);
        udf_comma_b     : in     vl_logic_vector(9 downto 0);
        udf_comma_mask  : in     vl_logic_vector(9 downto 0);
        uc_mode         : in     vl_logic;
        fc_mode         : in     vl_logic;
        pcie_mode       : in     vl_logic;
        rio_mode        : in     vl_logic;
        xge_mode        : in     vl_logic;
        ge_mode         : in     vl_logic;
        lsm_disable     : in     vl_logic;
        dec_bypass      : in     vl_logic;
        ctc_bypass      : in     vl_logic;
        ge_xmit         : in     vl_logic;
        ge_an_enable    : in     vl_logic;
        match1_d        : in     vl_logic_vector(9 downto 0);
        match2_d        : in     vl_logic_vector(9 downto 0);
        match3_d        : in     vl_logic_vector(9 downto 0);
        match4_d        : in     vl_logic_vector(9 downto 0);
        match2_en       : in     vl_logic;
        match4_en       : in     vl_logic;
        min_ipg_cnt     : in     vl_logic_vector(1 downto 0);
        high_mark       : in     vl_logic_vector(3 downto 0);
        low_mark        : in     vl_logic_vector(3 downto 0);
        cc_overrun      : out    vl_logic;
        cc_underrun     : out    vl_logic;
        pcie_det_done   : in     vl_logic;
        pcie_connect    : in     vl_logic;
        BISTRUN_A1      : in     vl_logic;
        BISTFC_A1       : in     vl_logic;
        BISTDONE_A1     : out    vl_logic;
        BISTF_A1        : out    vl_logic
    );
end pp_rx_top;
