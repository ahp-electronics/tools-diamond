library verilog;
use verilog.vl_types.all;
entity pcs_channel_top is
    generic(
        TIE_LO_STS      : integer := 0
    );
    port(
        sysclk          : in     vl_logic;
        sys_txrst_n     : in     vl_logic;
        sys_rxrst_n     : in     vl_logic;
        rxclk           : in     vl_logic;
        rxrst_n         : in     vl_logic;
        m_rxclk         : in     vl_logic;
        m_rxrst_n       : in     vl_logic;
        fb_rxclk        : in     vl_logic;
        fb_rxrst_n      : in     vl_logic;
        ff_tclk         : in     vl_logic;
        ff_rclk         : in     vl_logic;
        serdes_rxd      : in     vl_logic_vector(9 downto 0);
        sb_txd          : out    vl_logic_vector(9 downto 0);
        ff_txd          : in     vl_logic_vector(23 downto 0);
        fb_rxd          : out    vl_logic_vector(23 downto 0);
        x4_mode         : in     vl_logic;
        x2_mode         : in     vl_logic;
        mca_rxd_i       : in     vl_logic_vector(11 downto 0);
        mca_rxd_o       : out    vl_logic_vector(11 downto 0);
        t_detect_dni    : in     vl_logic;
        t_detect_upi    : in     vl_logic;
        t_detect_dno    : out    vl_logic;
        t_detect_upo    : out    vl_logic;
        align_status    : in     vl_logic;
        local_fault     : in     vl_logic_vector(8 downto 0);
        tx_slave        : in     vl_logic;
        rx_slave_x4     : in     vl_logic;
        rx_slave_x2     : in     vl_logic;
        idle_i          : in     vl_logic;
        a_count_i       : in     vl_logic_vector(4 downto 0);
        next_ifg_i      : in     vl_logic;
        code_sel_i      : in     vl_logic;
        seq_i           : in     vl_logic;
        idle_o          : out    vl_logic;
        a_count_o       : out    vl_logic_vector(4 downto 0);
        next_ifg_o      : out    vl_logic;
        code_sel_o      : out    vl_logic;
        seq_o           : out    vl_logic;
        cc_re_o         : out    vl_logic;
        cc_we_o         : out    vl_logic;
        cc_re_i         : in     vl_logic;
        cc_we_i         : in     vl_logic;
        fb_rxrst_i      : in     vl_logic;
        fb_rxrst_o      : out    vl_logic;
        fb_txrst_i      : in     vl_logic;
        fb_txrst_o      : out    vl_logic;
        ffc_signal_detect: in     vl_logic;
        ffc_enable_cgalign: in     vl_logic;
        ffc_fb_loopback : in     vl_logic;
        ffc_sb_inv_rx   : in     vl_logic;
        ffc_pcie_disable_tx: in     vl_logic;
        ffc_pcie_disable_rx: in     vl_logic;
        ls_sync_status  : out    vl_logic;
        ffs_cc_overrun  : out    vl_logic;
        ffs_cc_underrun : out    vl_logic;
        pcs_bypass      : in     vl_logic;
        pcs_mode        : in     vl_logic;
        fb_tx_mode      : in     vl_logic;
        fb_rx_mode      : in     vl_logic;
        xge_mode        : in     vl_logic;
        uc_mode         : in     vl_logic;
        pcie_mode       : in     vl_logic;
        rio_mode        : in     vl_logic;
        fc_mode         : in     vl_logic;
        lsm_disable     : in     vl_logic;
        udf_comma_a     : in     vl_logic_vector(9 downto 0);
        udf_comma_b     : in     vl_logic_vector(9 downto 0);
        udf_comma_mask  : in     vl_logic_vector(9 downto 0);
        match1_d        : in     vl_logic_vector(9 downto 0);
        match2_d        : in     vl_logic_vector(9 downto 0);
        match3_d        : in     vl_logic_vector(9 downto 0);
        match4_d        : in     vl_logic_vector(9 downto 0);
        match2_en       : in     vl_logic;
        match4_en       : in     vl_logic;
        min_ipg_cnt     : in     vl_logic_vector(1 downto 0);
        cc_hwm          : in     vl_logic_vector(3 downto 0);
        cc_lwm          : in     vl_logic_vector(3 downto 0);
        pcie_scram_select: in     vl_logic;
        prbs_select     : in     vl_logic;
        txcrc_swp       : in     vl_logic;
        txcrc_inv       : in     vl_logic;
        txcrc_swp_din   : in     vl_logic;
        txcrc_inv_din   : in     vl_logic;
        rxcrc_swp_din   : in     vl_logic;
        rxcrc_inv_din   : in     vl_logic;
        rxcrc_sopmk     : in     vl_logic_vector(8 downto 0);
        rxcrc_sopch_0   : in     vl_logic_vector(8 downto 0);
        rxcrc_sopch_1   : in     vl_logic_vector(8 downto 0);
        rxcrc_eopmk     : in     vl_logic_vector(8 downto 0);
        rxcrc_eopch_0   : in     vl_logic_vector(8 downto 0);
        rxcrc_eopch_1   : in     vl_logic_vector(8 downto 0);
        rxcrc_1ch       : in     vl_logic;
        rxcrc_swp_crc   : in     vl_logic;
        rxcrc_inv_crc   : in     vl_logic;
        rxcrc_swp_bytes : in     vl_logic;
        crc_initial     : in     vl_logic;
        crc_mode        : in     vl_logic_vector(1 downto 0);
        force_int       : in     vl_logic;
        rpwdnb          : out    vl_logic;
        tpwdnb          : out    vl_logic;
        rate_mode_rx    : out    vl_logic;
        rate_mode_tx    : out    vl_logic;
        rx_sdi_en       : out    vl_logic;
        tdrv_pre_en     : out    vl_logic;
        tdrv_pre_set    : out    vl_logic_vector(2 downto 0);
        rterm_tx        : out    vl_logic_vector(1 downto 0);
        tdrv_amp        : out    vl_logic_vector(1 downto 0);
        rterm_rx        : out    vl_logic_vector(1 downto 0);
        rcv_dcc_en      : out    vl_logic;
        req_en          : out    vl_logic;
        req_lvl_set     : out    vl_logic;
        rlol            : in     vl_logic;
        rlos_lo         : in     vl_logic;
        rlos_hi         : in     vl_logic;
        pcie_connect    : in     vl_logic;
        pcie_det_done   : in     vl_logic;
        sb_loopback     : out    vl_logic;
        rx_ch           : out    vl_logic;
        sonet_fbrx_mode : in     vl_logic;
        sonet_fbrx_wrst_n: in     vl_logic;
        sonet_fbrx_rrst_n: in     vl_logic;
        addro           : out    vl_logic_vector(7 downto 0);
        rdo             : out    vl_logic;
        wdatao          : out    vl_logic_vector(7 downto 0);
        wstbo           : out    vl_logic;
        rdatao          : out    vl_logic_vector(7 downto 0);
        into            : out    vl_logic;
        addri           : in     vl_logic_vector(7 downto 0);
        wdatai          : in     vl_logic_vector(7 downto 0);
        rdi             : in     vl_logic;
        wstbi           : in     vl_logic;
        rdatai          : in     vl_logic_vector(7 downto 0);
        inti            : in     vl_logic;
        int_cha_out     : out    vl_logic;
        cs_chif         : in     vl_logic;
        chif_rst_n      : in     vl_logic;
        bistrun_a1      : in     vl_logic;
        bistfc_a1       : in     vl_logic;
        bistdone_a1     : out    vl_logic_vector(1 downto 0);
        bistf_a1        : out    vl_logic_vector(1 downto 0);
        scan_mode       : in     vl_logic;
        scan_in_tx      : in     vl_logic;
        scan_in_rx      : in     vl_logic;
        scan_out_tx     : out    vl_logic;
        scan_out_rx     : out    vl_logic;
        char_td         : in     vl_logic_vector(9 downto 0);
        char_test_mode  : in     vl_logic_vector(2 downto 0)
    );
end pcs_channel_top;
