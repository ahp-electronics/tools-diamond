library verilog;
use verilog.vl_types.all;
entity FMCLK_TREE is
    port(
        A               : in     vl_logic;
        Z               : out    vl_logic
    );
end FMCLK_TREE;
