library verilog;
use verilog.vl_types.all;
entity ebr_polaritycntl is
    port(
        async_fuse      : in     vl_logic;
        f_grdis         : in     vl_logic;
        f_fifo_en       : in     vl_logic;
        gsrn            : in     vl_logic;
        gwe             : in     vl_logic;
        rsta            : in     vl_logic;
        f_prsta         : in     vl_logic;
        rstb            : in     vl_logic;
        f_prstb         : in     vl_logic;
        es_mode_rstn    : in     vl_logic;
        por_n           : in     vl_logic;
        cib_clka        : in     vl_logic;
        cib_clkb        : in     vl_logic;
        ebr_clkb        : in     vl_logic;
        f_mfg_clka      : in     vl_logic_vector(1 downto 0);
        f_mfg_clkb      : in     vl_logic_vector(1 downto 0);
        cea             : in     vl_logic;
        ceb             : in     vl_logic;
        oprcea          : in     vl_logic;
        oprceb          : in     vl_logic;
        w_ra            : in     vl_logic;
        f_pw_ra         : in     vl_logic;
        w_rb            : in     vl_logic;
        f_pw_rb         : in     vl_logic;
        cfg_cs          : in     vl_logic;
        csa             : in     vl_logic_vector(2 downto 0);
        f_pcsa          : in     vl_logic_vector(2 downto 0);
        csb             : in     vl_logic_vector(2 downto 0);
        f_pcsb          : in     vl_logic_vector(2 downto 0);
        es_mode         : in     vl_logic;
        f_rst_sync_dis  : in     vl_logic;
        async           : out    vl_logic;
        prsta           : out    vl_logic;
        prsta_del       : out    vl_logic;
        prsta_lookahead : out    vl_logic;
        prstb           : out    vl_logic;
        prstb_del       : out    vl_logic;
        prstb_lookahead : out    vl_logic;
        or_rstb         : out    vl_logic;
        ir_rsta         : out    vl_logic;
        ir_rstb         : out    vl_logic;
        pclka           : out    vl_logic;
        pclkb           : out    vl_logic;
        pcea            : out    vl_logic;
        pceb            : out    vl_logic;
        poprclka        : out    vl_logic;
        poprclkb        : out    vl_logic;
        poprcea         : out    vl_logic;
        poprceb         : out    vl_logic;
        porbuf          : out    vl_logic;
        pw_ra           : out    vl_logic;
        pw_rb           : out    vl_logic;
        pcsa            : out    vl_logic;
        pcsb            : out    vl_logic
    );
end ebr_polaritycntl;
