library verilog;
use verilog.vl_types.all;
entity e2bis_spare_gate is
    port(
        signal_in       : in     vl_logic
    );
end e2bis_spare_gate;
