-- $Header: //synplicity/map202003lat/mappers/cpld/lib/gen_mach/inc.vhd#1 $
@ER--HRMO:FRl8CkDRMoCC0sNFVsRHRDCVRFs#CkbsFOFDN5D0O0HC#RHbBvq]j6jj2vX
H
DLssN$ RQ 
 ;kR#CQ   38#0_oDFH4O_43ncN;DD
-

-----------------------------------------------------
R
CHM00Q$RhHBR#
R
oCCMs5HOMRR:HCM0o:Cs=c462
;R
sbF0
5R
:qRRRHM#_08DHFoOC_POs0F54M-RI8FMR0FjR2;
R
1:kRF00R#8F_Do_HOP0COFMs5-84RF0IMF2RjR2

;
R
CRM8Q;hBRN

sHOE00COkRsCpQe_hFBRVhRQB#RH
F
OlMbFCRM0e
BBRbRRF5s0
RRRRXRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR:R0FkR1RRap7_mBtQRR:='24';M
C8FROlMbFC;M0
F
OlMbFCRM0t
h7RbRRF5s0
RRRRXRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR:R0FkR1RRap7_mBtQRR:='2j';M
C8FROlMbFC;M0
F
OlMbFCRM0B_Bzq
77RbRRF5s0
RRRRqRRjRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR:RRHMR1RRap7_mBtQ;R
RRRRRARjRRRRRRRRRRRRRRRRRRRRRRRRRR:RRRMRHRRRR1_a7pQmtBR;
RRRRRhBQRRRRRRRRRRRRRRRRRRRRRRRRRRRR:HRRMRRRR71a_tpmQ
B;RRRRRjR1RRRRRRRRRRRRRRRRRRRRRRRRRRRRRR:RFRk0RaR17m_pt;QB
RRRRBRRmRzaRRRRRRRRRRRRRRRRRRRRRRRRRRR:R0FkR1RRap7_mBtQ2C;
MO8RFFlbM0CM;


#MHoNODRN$ssR:RRR8#0_oDFHPO_CFO0sM5R-84RF0IMFRRj2#;
HNoMDFROM_#04RR:#_08DHFoO#;
HNoMDFROM_#0jRR:#_08DHFoO
;
LHCoMz
S4e:RBuBRmR)av5quR>X=RMOF#40_2S;
zR.:tRh7uam)RuvqRR5X=O>RF0M#_;j2
RRRRRRRR:zdRzBB_7q7R)umaqRvuq5R5,j2RMOF#j0_,FROM_#041,R5,j2RsONsj$52
2;RRRRRRRRzRc:VRFsHMRHR04RF-RM4CRoMNCs0RC
RRRRRRRRRRRRRzRR.4_pRB:RBqz_7u7RmR)av5quRHq52O,RF0M#_Rj,OsNs$-5H4R2,125H,NROs5s$H;22
RRRRRRRR8CMRMoCC0sNC
;
CRM8pQe_h
B;
