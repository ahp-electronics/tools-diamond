library verilog;
use verilog.vl_types.all;
entity jtag_qual is
    port(
        isc_data_shift_iq: out    vl_logic;
        isc_addr_shift_iq: out    vl_logic;
        verify_id_iq    : out    vl_logic;
        idcode_pub_iq   : out    vl_logic;
        uidcode_pub_iq  : out    vl_logic;
        usercode_iq     : out    vl_logic;
        usercode_dryrun_iq: out    vl_logic;
        prog_dryrun_addr_iq: out    vl_logic;
        read_temp_iq    : out    vl_logic;
        idcode_prv_iq   : out    vl_logic;
        lsc_shift_password_iq: out    vl_logic;
        lsc_read_status_mq: out    vl_logic;
        lsc_read_status1_iq: out    vl_logic;
        lsc_read_mfg_status_mq: out    vl_logic;
        lsc_refresh_iq  : out    vl_logic;
        lsc_bitstream_burst_iq: out    vl_logic;
        lsc_i2ci_crbr_wt_iq: out    vl_logic;
        lsc_i2ci_txdr_wt_iq: out    vl_logic;
        lsc_i2ci_rxdr_rd_iq: out    vl_logic;
        lsc_i2ci_sr_rd_iq: out    vl_logic;
        lsc_read_pes_mq : out    vl_logic;
        lsc_device_ctrl_iq: out    vl_logic;
        lsc_prog_ctrl0_iq: out    vl_logic;
        lsc_read_ctrl0_iq: out    vl_logic;
        lsc_prog_ctrl1_iq: out    vl_logic;
        lsc_read_ctrl1_iq: out    vl_logic;
        lsc_reset_crc_iq: out    vl_logic;
        lsc_read_crc_iq : out    vl_logic;
        lsc_write_comp_dic_iq: out    vl_logic;
        lsc_read_comp_dic_mq: out    vl_logic;
        sf_prog_ucode_iq: out    vl_logic;
        sf_program_iq   : out    vl_logic;
        sf_read_iq      : out    vl_logic;
        sf_erase_iq     : out    vl_logic;
        sf_prog_done_iq : out    vl_logic;
        sf_erase_done_iq: out    vl_logic;
        sf_prog_sec_iq  : out    vl_logic;
        sf_init_addr_iq : out    vl_logic;
        sf_write_addr_iq: out    vl_logic;
        sf_prog_incr_rti_iq: out    vl_logic;
        sf_prog_incr_enc_iq: out    vl_logic;
        sf_prog_incr_cmp_iq: out    vl_logic;
        sf_prog_incr_cne_iq: out    vl_logic;
        sf_vfy_incr_rti_iq: out    vl_logic;
        sf_prog_sed_crc_iq: out    vl_logic;
        sf_read_sed_crc_iq: out    vl_logic;
        sf_write_bus_addr_iq: out    vl_logic;
        sf_pcs_write_iq : out    vl_logic;
        sf_pcs_read_iq  : out    vl_logic;
        sf_ebr_write_iq : out    vl_logic;
        sf_ebr_read_iq  : out    vl_logic;
        fl_prog_ucode_iq: out    vl_logic;
        fl_erase_iq     : out    vl_logic;
        fl_prog_done_iq : out    vl_logic;
        fl_prog_sec_iq  : out    vl_logic;
        fl_prog_secplus_iq: out    vl_logic;
        fl_init_addr_iq : out    vl_logic;
        fl_write_addr_iq: out    vl_logic;
        fl_prog_incr_nv_iq: out    vl_logic;
        fl_read_incr_nv_iq: out    vl_logic;
        fl_prog_password_iq: out    vl_logic;
        fl_read_password_iq: out    vl_logic;
        fl_prog_cipher_key0_iq: out    vl_logic;
        fl_read_cipher_key0_iq: out    vl_logic;
        fl_prog_cipher_key1_iq: out    vl_logic;
        fl_read_cipher_key1_iq: out    vl_logic;
        fl_prog_feature_iq: out    vl_logic;
        fl_read_feature_iq: out    vl_logic;
        fl_prog_feabits_iq: out    vl_logic;
        fl_read_feabits_iq: out    vl_logic;
        fl_init_addr_ufm_iq: out    vl_logic;
        fl_prog_tag_iq  : out    vl_logic;
        fl_erase_tag_iq : out    vl_logic;
        fl_read_tag_iq  : out    vl_logic;
        fl_prog_pes_mq  : out    vl_logic;
        fl_prog_trim0_mq: out    vl_logic;
        fl_prog_trim1_mq: out    vl_logic;
        fl_prog_mes_mq  : out    vl_logic;
        fl_prog_hes_mq  : out    vl_logic;
        fl_read_trim0_mq: out    vl_logic;
        fl_read_trim1_mq: out    vl_logic;
        fl_read_mes_mq  : out    vl_logic;
        fl_read_hes_mq  : out    vl_logic;
        fl_prog_csec_iq : out    vl_logic;
        fl_read_csec_iq : out    vl_logic;
        fl_prog_usec_iq : out    vl_logic;
        fl_read_usec_iq : out    vl_logic;
        fl_prog_authdone_iq: out    vl_logic;
        fl_prog_authmode_iq: out    vl_logic;
        fl_prog_aesfea_iq: out    vl_logic;
        fl_read_authmode_iq: out    vl_logic;
        fl_read_aesfea_iq: out    vl_logic;
        mfg_mtest_mq    : out    vl_logic;
        mfg_mtrim_mq    : out    vl_logic;
        mfg_mdata_mq    : out    vl_logic;
        mfg_bist_en_mq  : out    vl_logic;
        mfg_bist_status_mq: out    vl_logic;
        fl_prog_pubkey0_iq: out    vl_logic;
        fl_read_pubkey0_iq: out    vl_logic;
        fl_prog_pubkey1_iq: out    vl_logic;
        fl_read_pubkey1_iq: out    vl_logic;
        fl_prog_pubkey2_iq: out    vl_logic;
        fl_read_pubkey2_iq: out    vl_logic;
        fl_prog_pubkey3_iq: out    vl_logic;
        fl_read_pubkey3_iq: out    vl_logic;
        isc_enabled     : in     vl_logic;
        jaccess_sram    : in     vl_logic;
        jaccess_flash   : in     vl_logic;
        jaccess_tag     : in     vl_logic;
        jenable_tran    : in     vl_logic;
        ctrl_tran_edit  : in     vl_logic;
        mfg_en          : in     vl_logic;
        verify_id_i     : in     vl_logic;
        idcode_pub_i    : in     vl_logic;
        uidcode_pub_i   : in     vl_logic;
        usercode_i      : in     vl_logic;
        usercode_dryrun_i: in     vl_logic;
        prog_dryrun_addr_i: in     vl_logic;
        read_temp_i     : in     vl_logic;
        lsc_device_ctrl_i: in     vl_logic;
        lsc_shift_password_i: in     vl_logic;
        lsc_refresh_i   : in     vl_logic;
        lsc_bitstream_burst_i: in     vl_logic;
        lsc_i2ci_crbr_wt_i: in     vl_logic;
        lsc_i2ci_txdr_wt_i: in     vl_logic;
        lsc_i2ci_rxdr_rd_i: in     vl_logic;
        lsc_i2ci_sr_rd_i: in     vl_logic;
        idcode_prv_i    : in     vl_logic;
        isc_program_i   : in     vl_logic;
        isc_prog_ucode_i: in     vl_logic;
        isc_read_i      : in     vl_logic;
        isc_erase_i     : in     vl_logic;
        isc_prog_done_i : in     vl_logic;
        isc_erase_done_i: in     vl_logic;
        isc_prog_sec_i  : in     vl_logic;
        isc_prog_secplus_i: in     vl_logic;
        isc_data_shift_i: in     vl_logic;
        isc_addr_shift_i: in     vl_logic;
        lsc_init_addr_i : in     vl_logic;
        lsc_write_addr_i: in     vl_logic;
        lsc_prog_incr_rti_i: in     vl_logic;
        lsc_prog_incr_enc_i: in     vl_logic;
        lsc_prog_incr_cmp_i: in     vl_logic;
        lsc_prog_incr_cne_i: in     vl_logic;
        lsc_vfy_incr_rti_i: in     vl_logic;
        lsc_prog_ctrl0_i: in     vl_logic;
        lsc_read_ctrl0_i: in     vl_logic;
        lsc_prog_ctrl1_i: in     vl_logic;
        lsc_read_ctrl1_i: in     vl_logic;
        lsc_reset_crc_i : in     vl_logic;
        lsc_read_crc_i  : in     vl_logic;
        lsc_prog_sed_crc_i: in     vl_logic;
        lsc_read_sed_crc_i: in     vl_logic;
        lsc_prog_password_i: in     vl_logic;
        lsc_read_password_i: in     vl_logic;
        lsc_prog_cipher_key0_i: in     vl_logic;
        lsc_read_cipher_key0_i: in     vl_logic;
        lsc_prog_cipher_key1_i: in     vl_logic;
        lsc_read_cipher_key1_i: in     vl_logic;
        lsc_prog_feature_i: in     vl_logic;
        lsc_read_feature_i: in     vl_logic;
        lsc_prog_feabits_i: in     vl_logic;
        lsc_read_feabits_i: in     vl_logic;
        lsc_write_comp_dic_i: in     vl_logic;
        lsc_write_bus_addr_i: in     vl_logic;
        lsc_pcs_write_i : in     vl_logic;
        lsc_pcs_read_i  : in     vl_logic;
        lsc_ebr_write_i : in     vl_logic;
        lsc_ebr_read_i  : in     vl_logic;
        lsc_prog_incr_nv_i: in     vl_logic;
        lsc_read_incr_nv_i: in     vl_logic;
        lsc_init_addr_ufm_i: in     vl_logic;
        lsc_prog_tag_i  : in     vl_logic;
        lsc_erase_tag_i : in     vl_logic;
        lsc_read_tag_i  : in     vl_logic;
        lsc_prog_csec_i : in     vl_logic;
        lsc_read_csec_i : in     vl_logic;
        lsc_prog_usec_i : in     vl_logic;
        lsc_read_usec_i : in     vl_logic;
        lsc_prog_authdone_i: in     vl_logic;
        lsc_prog_authmode_i: in     vl_logic;
        lsc_prog_aesfea_i: in     vl_logic;
        lsc_read_authmode_i: in     vl_logic;
        lsc_read_aesfea_i: in     vl_logic;
        lsc_mtest_i     : in     vl_logic;
        lsc_mtrim_i     : in     vl_logic;
        lsc_mdata_i     : in     vl_logic;
        lsc_bist_en_i   : in     vl_logic;
        lsc_bist_status_i: in     vl_logic;
        lsc_read_status_m: in     vl_logic;
        lsc_read_mfg_status_m: in     vl_logic;
        lsc_read_status1_i: in     vl_logic;
        lsc_read_pes_m  : in     vl_logic;
        lsc_read_mes_m  : in     vl_logic;
        lsc_read_hes_m  : in     vl_logic;
        lsc_read_trim0_m: in     vl_logic;
        lsc_read_trim1_m: in     vl_logic;
        lsc_read_comp_dic_m: in     vl_logic;
        lsc_prog_pes_m  : in     vl_logic;
        lsc_prog_mes_m  : in     vl_logic;
        lsc_prog_hes_m  : in     vl_logic;
        lsc_prog_trim0_m: in     vl_logic;
        lsc_prog_trim1_m: in     vl_logic;
        lsc_prog_ecdsa_pubkey0_i: in     vl_logic;
        lsc_read_ecdsa_pubkey0_i: in     vl_logic;
        lsc_prog_ecdsa_pubkey1_i: in     vl_logic;
        lsc_read_ecdsa_pubkey1_i: in     vl_logic;
        lsc_prog_ecdsa_pubkey2_i: in     vl_logic;
        lsc_read_ecdsa_pubkey2_i: in     vl_logic;
        lsc_prog_ecdsa_pubkey3_i: in     vl_logic;
        lsc_read_ecdsa_pubkey3_i: in     vl_logic
    );
end jtag_qual;
