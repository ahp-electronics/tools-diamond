library verilog;
use verilog.vl_types.all;
entity sentry_flash is
    generic(
        CFG_ROWS        : integer := 272;
        UFM_ROWS        : integer := 64;
        TRIM_ROWS       : integer := 6;
        FEAT_ROWS       : integer := 6;
        COLUMNS         : integer := 1024;
        CFGFILE         : string  := "config.txt";
        UFMFILE         : string  := "ufm.txt";
        TRMFILE         : string  := "trim.txt";
        FEAFILE         : string  := "feat.txt"
    );
    port(
        fl_dout         : out    vl_logic_vector(63 downto 0);
        fl_ready        : out    vl_logic;
        fl_ready_por_n  : out    vl_logic;
        c_bl            : out    vl_logic_vector(3 downto 0);
        lastcol         : out    vl_logic_vector(3 downto 0);
        neg_edge_det    : out    vl_logic;
        well_active     : out    vl_logic;
        ready_vfy       : out    vl_logic;
        vwlp_active     : out    vl_logic;
        pumposc_mntr    : out    vl_logic;
        vpp_pos         : out    vl_logic;
        vpp_neg         : out    vl_logic;
        vread           : out    vl_logic;
        pos_mon         : out    vl_logic;
        well_pad        : out    vl_logic;
        l_row_cfg       : out    vl_logic;
        l_row_ufm       : out    vl_logic;
        vwlp_pad        : out    vl_logic;
        ufmrow_pad      : out    vl_logic;
        row             : in     vl_logic_vector(14 downto 0);
        ufm_row_sel_all : in     vl_logic;
        ufm_row_sel_none: in     vl_logic;
        cfg_row_sel_all : in     vl_logic;
        cfg_row_sel_none: in     vl_logic;
        trim_row_sel_all: in     vl_logic;
        trim_row_sel_none: in     vl_logic;
        feat_row_sel_all: in     vl_logic;
        feat_row_sel_none: in     vl_logic;
        era_ufm         : in     vl_logic;
        era_cfg         : in     vl_logic;
        era_trim        : in     vl_logic;
        era_feat        : in     vl_logic;
        prg_ufm         : in     vl_logic;
        prg_cfg         : in     vl_logic;
        prg_tf          : in     vl_logic;
        read_ufm        : in     vl_logic;
        read_cfg        : in     vl_logic;
        read_tf         : in     vl_logic;
        erase_setup     : in     vl_logic;
        erapdis         : in     vl_logic;
        erase_pulse     : in     vl_logic;
        pwtc_well       : in     vl_logic;
        prg_pulse       : in     vl_logic_vector(3 downto 0);
        prog_disch      : in     vl_logic;
        prg_pwtc        : in     vl_logic;
        en_vreg_mon     : in     vl_logic;
        era_ver         : in     vl_logic;
        scp             : in     vl_logic;
        softprg         : in     vl_logic;
        verify          : in     vl_logic;
        flash_en        : in     vl_logic;
        reg_enable      : in     vl_logic;
        subrow_mvena_ufm: in     vl_logic;
        subrow_mvenall_ufm: in     vl_logic;
        subrow_hvena_ufm: in     vl_logic;
        subrow_hvenall_ufm: in     vl_logic;
        subrow_mvena_cfg: in     vl_logic;
        subrow_mvenall_cfg: in     vl_logic;
        subrow_hvena_cfg: in     vl_logic;
        subrow_hvenall_cfg: in     vl_logic;
        subrow_mvena_tf : in     vl_logic;
        subrow_hvena_tf : in     vl_logic;
        sa_enall        : in     vl_logic;
        sa_ena          : in     vl_logic;
        prgdrv_enall    : in     vl_logic;
        prgdrv_ena      : in     vl_logic;
        col_shift       : in     vl_logic;
        colstart        : in     vl_logic_vector(3 downto 0);
        col_rst         : in     vl_logic;
        readpart        : in     vl_logic_vector(3 downto 0);
        wor_eval        : in     vl_logic;
        wand_eval       : in     vl_logic;
        capture_dout    : in     vl_logic;
        src_clamp       : in     vl_logic;
        scpv            : in     vl_logic;
        drain_ctrl      : in     vl_logic;
        ppt_en          : in     vl_logic;
        ppt_pset        : in     vl_logic;
        ppt_rowsel      : in     vl_logic;
        sel_6p5v        : in     vl_logic;
        prestep_in_neg  : in     vl_logic_vector(2 downto 0);
        step_in_neg     : in     vl_logic_vector(2 downto 0);
        margin_in       : in     vl_logic;
        fl_ready_rst    : in     vl_logic;
        por_init_n      : in     vl_logic;
        vccaux          : in     vl_logic;
        mfg_negpumpoff  : in     vl_logic;
        mfg_vread0_n    : in     vl_logic;
        mfg_vpp_n       : in     vl_logic;
        mfg_well_obs    : in     vl_logic;
        mfg_vpos_mon    : in     vl_logic;
        mfg_vread_mon   : in     vl_logic;
        mfg_vwlp_mon    : in     vl_logic;
        vpos_trim       : in     vl_logic_vector(4 downto 0);
        vpp_trim        : in     vl_logic_vector(3 downto 0);
        vread_trim      : in     vl_logic_vector(3 downto 0);
        vreg_trim       : in     vl_logic_vector(2 downto 0);
        neg_pump_sel    : in     vl_logic;
        trim_src_res    : in     vl_logic_vector(1 downto 0);
        shared_iref_bias: in     vl_logic;
        i10ua_4vref     : in     vl_logic;
        mfg_vwlp_obs    : in     vl_logic;
        mfg_ufmwl_obs   : in     vl_logic;
        mfg_fl_spare3   : in     vl_logic;
        mfg_fl_spare4   : in     vl_logic;
        mfg_margin      : in     vl_logic;
        mfg_pumposc_oe  : in     vl_logic
    );
end sentry_flash;
