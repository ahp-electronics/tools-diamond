library verilog;
use verilog.vl_types.all;
entity pcs_quad_buffers is
    port(
        cyawstn         : in     vl_logic;
        tri_ion         : in     vl_logic;
        sciaddr         : in     vl_logic_vector(5 downto 0);
        scienaux        : in     vl_logic;
        sciench0        : in     vl_logic;
        sciench1        : in     vl_logic;
        sciench2        : in     vl_logic;
        sciench3        : in     vl_logic;
        scird           : in     vl_logic;
        sciselaux       : in     vl_logic;
        sciselch0       : in     vl_logic;
        sciselch1       : in     vl_logic;
        sciselch2       : in     vl_logic;
        sciselch3       : in     vl_logic;
        sciwdata        : in     vl_logic_vector(7 downto 0);
        sciwstn         : in     vl_logic;
        scienaux_b      : out    vl_logic;
        sciench0_b      : out    vl_logic;
        sciench1_b      : out    vl_logic;
        sciench2_b      : out    vl_logic;
        sciench3_b      : out    vl_logic;
        sciselaux_b     : out    vl_logic;
        sciselch0_b     : out    vl_logic;
        sciselch1_b     : out    vl_logic;
        sciselch2_b     : out    vl_logic;
        sciselch3_b     : out    vl_logic;
        scirdata        : out    vl_logic_vector(7 downto 0);
        sciint          : out    vl_logic;
        sci_resetn32    : out    vl_logic;
        sci_ion_dl32    : out    vl_logic;
        sci_wstb32      : out    vl_logic;
        sci_rd32        : out    vl_logic;
        sci_addr32      : out    vl_logic_vector(5 downto 0);
        sci_wdata32     : out    vl_logic_vector(7 downto 0);
        sci_rdata32     : in     vl_logic_vector(7 downto 0);
        sci_int32       : in     vl_logic;
        sci_resetn10    : out    vl_logic;
        sci_ion_dl10    : out    vl_logic;
        sci_wstb10      : out    vl_logic;
        sci_rd10        : out    vl_logic;
        sci_addr10      : out    vl_logic_vector(5 downto 0);
        sci_wdata10     : out    vl_logic_vector(7 downto 0);
        sci_rdata10     : in     vl_logic_vector(7 downto 0);
        sci_int10       : in     vl_logic;
        sci_resetnaux   : out    vl_logic;
        sci_ion_dlaux   : out    vl_logic;
        sci_wstbaux     : out    vl_logic;
        sci_rdaux       : out    vl_logic;
        sci_addraux     : out    vl_logic_vector(5 downto 0);
        sci_wdataaux    : out    vl_logic_vector(7 downto 0);
        sci_rdataaux    : in     vl_logic_vector(7 downto 0);
        sci_intaux      : in     vl_logic;
        tri_ion_reset   : out    vl_logic
    );
end pcs_quad_buffers;
