//
// Functional Coverage package
//

package mti_fcover;
    typedef enum {SYM = 1, BIN = 2, OCT = 8, DEC = 10, HEX = 16} mtiRadixKind;
endpackage
