-- $Header: //synplicity/map202003lat/mappers/lattice/lib/gen_lava1/cmp_lt.vhd#1 $
@ER--O_lbDD0
HNLssQ$R ;  
Ck#R Q  03#8F_Do_HO4c4n3DND;C

M00H$vRBua_pR
H#
MoCCOsH58IH0RE:HCM0o:Cs=d4.2
;
b0Fs5q

,:ARRRHM#_08DHFoOC_POs0F58IH04E-RI8FMR0Fj
2;
Rpa:kRF00R#8F_Do
HO

2;
8CMRuBv_;pa
s
NO0EHCkO0spCRev_Bua_pRRFVB_vupHaR#O

FFlbM0CMRzBB_Aqt
RRRb0Fs5R
RRRRRqRjRRRRRRRRRRRRRRRRRRRRRRRRRR:RRRMRHRRRR1_a7pQmtBR;
RRRRRRAjRRRRRRRRRRRRRRRRRRRRRRRRRRRR:HRRMRRRR71a_tpmQ
B;RRRRRQRBhRRRRRRRRRRRRRRRRRRRRRRRRRRRRR:RHRMRRaR17m_pt;QB
RRRRBRRmRzaRRRRRRRRRRRRRRRRRRRRRRRRRRR:R0FkR1RRap7_mBtQ2C;
MO8RFFlbM0CM;O

FFlbM0CMRBeB
RRRb0Fs5R
RRRRRXRRRRRRRRRRRRRRRRRRRRRRRRRRRR:RRRkRF0RRR1_a7pQmtB=R:R''j2C;
MO8RFFlbM0CM;O

FFlbM0CMReQh
RRRb0Fs5R
RRRRRQRjRRRRRRRRRRRRRRRRRRRRRRRRRR:RRRMRHRRRR1_a7pQmtBR;
RRRRRRmRRRRRRRRRRRRRRRRRRRRRRRRRRRRR:FRRkR0RR71a_tpmQ;B2
8CMRlOFbCFMM
0;
H
#oDMNRsONsR$RR#:R0D8_FOoH_OPC05FsR8IH04E-RI8FMR0Fj;R2
o#HMRNDO#FM0R_j:0R#8F_Do;HO
C
Lo
HMS:z4RBeBR)umaqRvuX5R=F>OM_#0j;R2
.Sz:BRBzt_qAmRu)vaRqRu5q>j=q25j,jRA=5>AjR2,B=Qh>MOF#j0_,mRBz>a=OsNs$25jR
2;S:zdRsVFRHHRMRR40IFRHE80-o4RCsMCN
0CSdSz_:p4RzBB_AqtR)umaqRvuq5Rjq=>5,H2R=Aj>HA52B,RQ>h=OsNs$-5H4R2,Bamz=N>Os5s$H22R;C
SMo8RCsMCN;0C
cSz:hRQemRu)vaRq5uRQ>j=RsONsI$5HE80R2-4,=Rm>2pa;C

Mp8Rev_Bua_p;



