library verilog;
use verilog.vl_types.all;
entity bsctl8_1 is
    port(
        TDO             : out    vl_logic;
        TDOE            : out    vl_logic;
        TDOEN           : out    vl_logic;
        PRGM_JTAG       : out    vl_logic;
        RD_CFG_JTAG     : out    vl_logic;
        TDI_JTAG        : out    vl_logic;
        ENTCK_JTAG      : out    vl_logic;
        JTAG_MODE       : out    vl_logic;
        BS_MODE         : out    vl_logic;
        INTEST          : out    vl_logic;
        HIGHZ           : out    vl_logic;
        SHBSRN          : out    vl_logic;
        CPTBSR          : out    vl_logic;
        UPDTBSR         : out    vl_logic;
        TRESET          : out    vl_logic;
        PSRSFTN         : out    vl_logic;
        PSRCAP          : out    vl_logic;
        TDI1_LASB       : out    vl_logic;
        TDI1_RASB       : out    vl_logic;
        SHDR            : out    vl_logic;
        CPTDR           : out    vl_logic;
        UPDTDR          : out    vl_logic;
        RUNTST          : out    vl_logic;
        DOBIST_LASB     : out    vl_logic;
        DOBIST_RASB     : out    vl_logic;
        PSRENABLE1      : out    vl_logic;
        PSRENABLE2      : out    vl_logic;
        PSRENABLE3      : out    vl_logic;
        SCANENABLE      : out    vl_logic_vector(16 downto 1);
        JRSTN           : out    vl_logic;
        JTCK            : out    vl_logic;
        JTDI            : out    vl_logic;
        JSHIFT          : out    vl_logic;
        JUPDATE         : out    vl_logic;
        JCE             : out    vl_logic_vector(8 downto 1);
        JRTI            : out    vl_logic_vector(8 downto 1);
        TCK             : in     vl_logic;
        TCKD            : in     vl_logic;
        TMS             : in     vl_logic;
        TDI             : in     vl_logic;
        BSRSO           : in     vl_logic;
        PIN_TSN         : in     vl_logic;
        SO_BIST_LASB    : in     vl_logic;
        SO_BIST_RASB    : in     vl_logic;
        VENDORID        : in     vl_logic_vector(31 downto 0);
        MC1_USERBIT     : in     vl_logic_vector(31 downto 0);
        CHIPID          : in     vl_logic_vector(7 downto 0);
        CFGDOUTN        : in     vl_logic;
        RDBK_DATA       : in     vl_logic;
        RDBK_TDO_EN     : in     vl_logic;
        PAD_DONE        : in     vl_logic;
        PSROUT1         : in     vl_logic;
        PSROUT2         : in     vl_logic;
        PSROUT3         : in     vl_logic;
        JTDO            : in     vl_logic_vector(8 downto 1);
        SCANOUT         : in     vl_logic_vector(16 downto 9);
        TS_ALL          : in     vl_logic;
        MC1_SCAN        : in     vl_logic_vector(8 downto 1);
        MC1_EN_SPI_N    : in     vl_logic;
        USR_TDO         : in     vl_logic;
        MC1_USR_TDO     : in     vl_logic
    );
end bsctl8_1;
