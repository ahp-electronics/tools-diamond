library verilog;
use verilog.vl_types.all;
entity X151T001 is
    port(
        VDDA            : inout  vl_logic;
        VSSA            : inout  vl_logic;
        VDD             : inout  vl_logic;
        VSS             : inout  vl_logic;
        DVSS            : inout  vl_logic;
        HSEL            : in     vl_logic;
        BITCLK          : in     vl_logic;
        PD              : in     vl_logic;
        PDBIAS          : in     vl_logic;
        LB_EN           : in     vl_logic;
        ENP_DESER       : in     vl_logic;
        PDCKG           : in     vl_logic;
        HS_16BIT_EN     : in     vl_logic;
        TX_RCAL         : in     vl_logic;
        RX_RCAL         : in     vl_logic_vector(1 downto 0);
        DP0             : inout  vl_logic;
        DN0             : inout  vl_logic;
        D0_DTXLPP       : in     vl_logic;
        D0_DTXLPN       : in     vl_logic;
        D0_TXLPEN       : in     vl_logic;
        D0_DRXLPP       : out    vl_logic;
        D0_DRXLPN       : out    vl_logic;
        D0_RXLPEN       : in     vl_logic;
        D0_DCDP         : out    vl_logic;
        D0_DCDN         : out    vl_logic;
        D0_CDEN         : in     vl_logic;
        D0_TXHSPD       : in     vl_logic;
        D0_TXHSEN       : in     vl_logic;
        D0_HSTX_DATA    : in     vl_logic_vector(15 downto 0);
        D0_HS_SER_EN    : in     vl_logic;
        D0_RXHSEN       : in     vl_logic;
        D0_HS_DESER_EN  : in     vl_logic;
        D0_HSRX_DATA    : out    vl_logic_vector(15 downto 0);
        D0_HS_BYTE_CLKD : out    vl_logic;
        D0_SYNC         : out    vl_logic;
        D0_ERRSYNC      : out    vl_logic;
        D0_NOSYNC       : out    vl_logic;
        D0_DRXHS        : out    vl_logic;
        D0_HS_BYTE_CLKS : out    vl_logic;
        DP1             : inout  vl_logic;
        DN1             : inout  vl_logic;
        D1_DTXLPP       : in     vl_logic;
        D1_DTXLPN       : in     vl_logic;
        D1_TXLPEN       : in     vl_logic;
        D1_DRXLPP       : out    vl_logic;
        D1_DRXLPN       : out    vl_logic;
        D1_RXLPEN       : in     vl_logic;
        D1_DCDP         : out    vl_logic;
        D1_DCDN         : out    vl_logic;
        D1_CDEN         : in     vl_logic;
        D1_TXHSPD       : in     vl_logic;
        D1_TXHSEN       : in     vl_logic;
        D1_HSTX_DATA    : in     vl_logic_vector(15 downto 0);
        D1_HS_SER_EN    : in     vl_logic;
        D1_RXHSEN       : in     vl_logic;
        D1_HS_DESER_EN  : in     vl_logic;
        D1_HSRX_DATA    : out    vl_logic_vector(15 downto 0);
        D1_SYNC         : out    vl_logic;
        D1_ERRSYNC      : out    vl_logic;
        D1_NOSYNC       : out    vl_logic;
        D1_DRXHS        : out    vl_logic;
        DP2             : inout  vl_logic;
        DN2             : inout  vl_logic;
        D2_DTXLPP       : in     vl_logic;
        D2_DTXLPN       : in     vl_logic;
        D2_TXLPEN       : in     vl_logic;
        D2_DRXLPP       : out    vl_logic;
        D2_DRXLPN       : out    vl_logic;
        D2_RXLPEN       : in     vl_logic;
        D2_DCDP         : out    vl_logic;
        D2_DCDN         : out    vl_logic;
        D2_CDEN         : in     vl_logic;
        D2_TXHSPD       : in     vl_logic;
        D2_TXHSEN       : in     vl_logic;
        D2_HSTX_DATA    : in     vl_logic_vector(15 downto 0);
        D2_HS_SER_EN    : in     vl_logic;
        D2_RXHSEN       : in     vl_logic;
        D2_HS_DESER_EN  : in     vl_logic;
        D2_HSRX_DATA    : out    vl_logic_vector(15 downto 0);
        D2_SYNC         : out    vl_logic;
        D2_ERRSYNC      : out    vl_logic;
        D2_NOSYNC       : out    vl_logic;
        D2_DRXHS        : out    vl_logic;
        DP3             : inout  vl_logic;
        DN3             : inout  vl_logic;
        D3_DTXLPP       : in     vl_logic;
        D3_DTXLPN       : in     vl_logic;
        D3_TXLPEN       : in     vl_logic;
        D3_DRXLPP       : out    vl_logic;
        D3_DRXLPN       : out    vl_logic;
        D3_RXLPEN       : in     vl_logic;
        D3_DCDP         : out    vl_logic;
        D3_DCDN         : out    vl_logic;
        D3_CDEN         : in     vl_logic;
        D3_TXHSPD       : in     vl_logic;
        D3_TXHSEN       : in     vl_logic;
        D3_HSTX_DATA    : in     vl_logic_vector(15 downto 0);
        D3_HS_SER_EN    : in     vl_logic;
        D3_RXHSEN       : in     vl_logic;
        D3_HS_DESER_EN  : in     vl_logic;
        D3_HSRX_DATA    : out    vl_logic_vector(15 downto 0);
        D3_SYNC         : out    vl_logic;
        D3_ERRSYNC      : out    vl_logic;
        D3_NOSYNC       : out    vl_logic;
        D3_DRXHS        : out    vl_logic;
        CKP             : inout  vl_logic;
        CKN             : inout  vl_logic;
        CLK_DTXLPP      : in     vl_logic;
        CLK_DTXLPN      : in     vl_logic;
        CLK_TXLPEN      : in     vl_logic;
        CLK_DRXLPP      : out    vl_logic;
        CLK_DRXLPN      : out    vl_logic;
        CLK_RXLPEN      : in     vl_logic;
        CLK_DCDN        : out    vl_logic;
        CLK_CDEN        : in     vl_logic;
        CLK_TXHSPD      : in     vl_logic;
        CLK_TXHSEN      : in     vl_logic;
        CLK_TXHSGATE    : in     vl_logic;
        CLK_RXHSEN      : in     vl_logic;
        CLK_HS_BYTE     : out    vl_logic;
        CLK_DRXHS       : out    vl_logic
    );
end X151T001;
