library verilog;
use verilog.vl_types.all;
entity config_cntl is
    port(
        tdo             : out    vl_logic;
        jshift          : out    vl_logic;
        jtdi            : out    vl_logic;
        jce             : out    vl_logic_vector(2 downto 1);
        por             : out    vl_logic;
        por_sec         : out    vl_logic;
        por_trim        : out    vl_logic;
        por_jtag        : out    vl_logic;
        scan_en_out     : out    vl_logic;
        scan_mode       : out    vl_logic;
        cfg_addr_por_n  : out    vl_logic;
        cfg_data_por_n  : out    vl_logic;
        sram_ppt_addr   : out    vl_logic_vector(3 downto 0);
        gsrn            : out    vl_logic;
        wb_dat_o        : out    vl_logic_vector(7 downto 0);
        scan_in         : out    vl_logic_vector(7 downto 0);
        tms             : in     vl_logic;
        tdi             : in     vl_logic;
        tdo_in          : in     vl_logic;
        programn_pin    : in     vl_logic;
        sf_ppt_addr     : in     vl_logic_vector(3 downto 0);
        isptcy_shcap    : in     vl_logic;
        isptcy_tdi      : in     vl_logic;
        isptcy_ener1    : in     vl_logic;
        isptcy_ener2    : in     vl_logic;
        iscan_en        : in     vl_logic_vector(7 downto 0);
        jtdo            : in     vl_logic_vector(2 downto 1);
        sed_frcerr      : in     vl_logic;
        pfsafe          : in     vl_logic;
        pwrup_pur_n     : in     vl_logic;
        cfg_osc         : in     vl_logic;
        smclk           : in     vl_logic;
        gsrn_sync_clk   : in     vl_logic;
        gsrn_out        : in     vl_logic;
        gsrn_sync       : in     vl_logic;
        mc1_scan_test_en: in     vl_logic_vector(3 downto 0);
        wb_dat_o_sci    : in     vl_logic_vector(7 downto 0);
        scan_out        : in     vl_logic_vector(7 downto 0);
        isc_exec_d      : in     vl_logic;
        wb_adr_i        : in     vl_logic_vector(7 downto 0);
        wb_cyc_i        : in     vl_logic;
        wb_we_i         : in     vl_logic;
        wb_clk_i        : in     vl_logic;
        cib_i2c_scl_i   : in     vl_logic;
        cib_i2c_sda_i   : in     vl_logic
    );
end config_cntl;
