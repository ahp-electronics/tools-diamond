library verilog;
use verilog.vl_types.all;
entity pcs_channel_top is
    port(
        bist_rx_data_sel: in     vl_logic;
        bistfc_a1       : in     vl_logic;
        bistrun_a1      : in     vl_logic;
        char_mode       : in     vl_logic;
        char_test_data  : in     vl_logic_vector(9 downto 0);
        char_test_mode  : in     vl_logic;
        ebrd_clk        : in     vl_logic;
        fb_clk          : in     vl_logic;
        fc_mode         : in     vl_logic;
        ff_ebrd_clk     : in     vl_logic;
        ff_rx_clk_sel   : in     vl_logic_vector(2 downto 0);
        ff_rxi_clk      : in     vl_logic;
        ff_tx_d         : in     vl_logic_vector(23 downto 0);
        ff_txi_clk      : in     vl_logic;
        ffc_ei_en       : in     vl_logic;
        ffc_enable_cgalign: in     vl_logic;
        ffc_fb_loopback : in     vl_logic;
        ffc_lane_rx_rst : in     vl_logic;
        ffc_lane_tx_rst : in     vl_logic;
        ffc_pcie_ct     : in     vl_logic;
        ffc_pfifo_clr   : in     vl_logic;
        ffc_rxpwdnb     : in     vl_logic;
        ffc_sb_inv_rx   : in     vl_logic;
        ffc_sb_pfifo_lp : in     vl_logic;
        ffc_signal_detect: in     vl_logic;
        ffc_txpwdnb     : in     vl_logic;
        ffr_clk         : in     vl_logic;
        fft_clk         : in     vl_logic;
        fmbist_data     : in     vl_logic_vector(9 downto 0);
        force_int       : in     vl_logic;
        ion_delay       : in     vl_logic;
        lane_rx_rst     : in     vl_logic;
        lane_tx_rst     : in     vl_logic;
        mc1_chif_ctl    : in     vl_logic_vector(103 downto 0);
        pcie_connect    : in     vl_logic;
        pcie_det_done   : in     vl_logic;
        pcie_mode       : in     vl_logic;
        pcs_addri       : in     vl_logic_vector(5 downto 0);
        pcs_ctl_10_qd_09: in     vl_logic_vector(7 downto 0);
        pcs_ctl_11_qd_0a: in     vl_logic_vector(7 downto 0);
        pcs_ctl_12_qd_0b: in     vl_logic_vector(7 downto 0);
        pcs_ctl_13_qd_0c: in     vl_logic_vector(7 downto 0);
        pcs_ctl_3_qd_02 : in     vl_logic_vector(7 downto 0);
        pcs_ctl_4_qd_03 : in     vl_logic_vector(7 downto 0);
        pcs_ctl_5_qd_04 : in     vl_logic_vector(7 downto 0);
        pcs_ctl_6_qd_05 : in     vl_logic_vector(7 downto 0);
        pcs_ctl_7_qd_06 : in     vl_logic_vector(7 downto 0);
        pcs_ctl_8_qd_07 : in     vl_logic_vector(7 downto 0);
        pcs_ctl_9_qd_08 : in     vl_logic_vector(7 downto 0);
        pcs_inti        : in     vl_logic;
        pcs_rdatai      : in     vl_logic_vector(7 downto 0);
        pcs_rdi         : in     vl_logic;
        pcs_wdatai      : in     vl_logic_vector(7 downto 0);
        pcs_wstbi       : in     vl_logic;
        plol            : in     vl_logic;
        quad_reset_all  : in     vl_logic;
        quad_reset_all_n: in     vl_logic;
        rio_mode        : in     vl_logic;
        rlol            : in     vl_logic;
        rlos_hi         : in     vl_logic;
        rlos_lo         : in     vl_logic;
        rlos_com        : out    vl_logic;
        rst_ebrd_clk_n  : in     vl_logic;
        rst_fb_clk_n    : in     vl_logic;
        rst_rx_clk_n    : in     vl_logic;
        rst_tx_clk_n    : in     vl_logic;
        rx_clk          : in     vl_logic;
        sci_resetn      : in     vl_logic;
        sciench         : in     vl_logic;
        sciselch        : in     vl_logic;
        sd_rx_clk       : in     vl_logic;
        sd_tx_clk       : in     vl_logic;
        sel_sd_rx_clk   : in     vl_logic;
        ser_sts_2_ch_27 : in     vl_logic_vector(7 downto 0);
        ser_sts_3_ch_28 : in     vl_logic_vector(7 downto 0);
        ser_sts_4_ch_29 : in     vl_logic_vector(7 downto 0);
        ser_sts_6_ch_2b : in     vl_logic_vector(7 downto 0);
        ser_sts_7_ch_2c : in     vl_logic_vector(7 downto 0);
        serdes_rxd      : in     vl_logic_vector(9 downto 0);
        test_clk        : in     vl_logic;
        tx_clk          : in     vl_logic;
        uc_mode         : in     vl_logic;
        xge_mode        : in     vl_logic;
        bistdone_a1     : out    vl_logic_vector(1 downto 0);
        bistf_a1        : out    vl_logic_vector(1 downto 0);
        ctie_low        : out    vl_logic;
        ebrd_clk_o      : out    vl_logic;
        fb_clk_o        : out    vl_logic;
        ff_rx_d         : out    vl_logic_vector(23 downto 0);
        ff_rx_f_clk     : out    vl_logic;
        ff_rx_h_clk     : out    vl_logic;
        ff_rx_q_clk     : out    vl_logic;
        ffr_clk_o       : out    vl_logic;
        ffs_cc_overrun  : out    vl_logic;
        ffs_cc_underrun : out    vl_logic;
        ffs_ls_sync_status: out    vl_logic;
        ffs_rxfbfifo_error: out    vl_logic;
        ffs_txfbfifo_error: out    vl_logic;
        fft_clk_o       : out    vl_logic;
        int_cha_out     : out    vl_logic;
        pcs_addro       : out    vl_logic_vector(5 downto 0);
        pcs_into        : out    vl_logic;
        pcs_rdatao      : out    vl_logic_vector(7 downto 0);
        pcs_rdo         : out    vl_logic;
        pcs_wdatao      : out    vl_logic_vector(7 downto 0);
        pcs_wstbo       : out    vl_logic;
        rst_ebrd_clk_n_o: out    vl_logic;
        rst_fb_clk_n_o  : out    vl_logic;
        rst_rx_clk_n_o  : out    vl_logic;
        rst_tx_clk_n_o  : out    vl_logic;
        rx_ch           : out    vl_logic;
        rx_clk_o        : out    vl_logic;
        sb_txd          : out    vl_logic_vector(9 downto 0);
        ser_ctl_1_ch_07 : out    vl_logic_vector(7 downto 0);
        ser_ctl_2_ch_08 : out    vl_logic_vector(7 downto 0);
        ser_ctl_3_ch_09 : out    vl_logic_vector(7 downto 0);
        ser_ctl_4_ch_0a : out    vl_logic_vector(7 downto 0);
        ser_ctl_5_ch_0b : out    vl_logic_vector(7 downto 0);
        tobist_data     : out    vl_logic_vector(9 downto 0);
        tsd_pcie_det_ct : out    vl_logic;
        tsd_pcie_ei_en  : out    vl_logic;
        tx_clk_o        : out    vl_logic
    );
end pcs_channel_top;
