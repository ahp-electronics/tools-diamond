library verilog;
use verilog.vl_types.all;
entity datap_unit is
    generic(
        COMP_DIC_LENGTH : integer := 16;
      --CR_SEED         : integer type with unrepresentable value!
        AES_MODE        : integer := 1
      --UDS_PADDING_BITS: integer type with unrepresentable value!
    );
    port(
        njtag_run       : out    vl_logic;
        nj_dat_ren      : out    vl_logic;
        nj_dat_wen      : out    vl_logic;
        njtag_din       : out    vl_logic_vector(7 downto 0);
        decompress_njtag_en: out    vl_logic;
        dec_load        : out    vl_logic;
        rfifo_re        : out    vl_logic;
        wfifo_we        : out    vl_logic;
        wfifo_din       : out    vl_logic_vector(7 downto 0);
        decompress_1byte: out    vl_logic;
        decompress_8byte: out    vl_logic;
        decompress_out  : out    vl_logic_vector(63 downto 0);
        decrypt_burst   : out    vl_logic;
        decrypt_out     : out    vl_logic_vector(7 downto 0);
        dp_dsr_8byte_cmp: out    vl_logic;
        dp_dsr_1byte_cmp: out    vl_logic;
        dp_dsr_1byte_enc: out    vl_logic;
        cfg_crc         : out    vl_logic_vector(15 downto 0);
        njm_crc_err     : out    vl_logic;
        sdm_run         : out    vl_logic;
        dec_init_done   : out    vl_logic;
        auth_init_done  : out    vl_logic;
        hse_clk         : in     vl_logic;
        hse_reset       : out    vl_logic;
        hse_enc_enable  : out    vl_logic;
        hse_cfg_active  : out    vl_logic;
        hse_cfg_noise   : out    vl_logic;
        hse_ac_alg_sel  : out    vl_logic_vector(1 downto 0);
        hse_data_in     : out    vl_logic_vector(7 downto 0);
        hse_write_en    : out    vl_logic;
        hse_last_byte   : out    vl_logic;
        auth_en         : out    vl_logic;
        auth_fail       : out    vl_logic;
        auth_done       : out    vl_logic;
        auth_time_out   : out    vl_logic;
        auth_setup_fail : out    vl_logic;
        auth_bs_err     : out    vl_logic;
        key_rst_sync    : out    vl_logic;
        key_shift_en    : out    vl_logic;
        hse_trn_dat     : out    vl_logic_vector(127 downto 0);
        hse_uds_in      : out    vl_logic_vector(255 downto 0);
        por             : in     vl_logic;
        por_sec         : in     vl_logic;
        smclk           : in     vl_logic;
        scan_mode       : in     vl_logic;
        isc_rst_sync    : in     vl_logic;
        sed_en_adv      : in     vl_logic;
        sed_active      : in     vl_logic;
        njtag_slv_en    : in     vl_logic;
        njfsm_hold      : in     vl_logic;
        jtag_active_smsync: in     vl_logic;
        ShiftDR         : in     vl_logic;
        isc_data_shift_iqual: in     vl_logic;
        lsc_prog_incr_rti_iqual: in     vl_logic;
        lsc_prog_incr_enc_iqual: in     vl_logic;
        lsc_prog_incr_cne_iqual: in     vl_logic;
        lsc_prog_incr_cmp_iqual: in     vl_logic;
        lsc_bitstream_burst_iq: in     vl_logic;
        njtag_active    : in     vl_logic;
        njtag_cmd       : in     vl_logic;
        njtag_infa      : in     vl_logic;
        njshf_dat0      : in     vl_logic;
        njshf_dat       : in     vl_logic;
        njshf_crc       : in     vl_logic;
        njshf_dum       : in     vl_logic;
        njbse_rxcmd     : in     vl_logic;
        njbse_rxdec     : in     vl_logic;
        isc_data_shift_cqual: in     vl_logic;
        lsc_prog_incr_rti_cqual: in     vl_logic;
        lsc_prog_incr_enc_cqual: in     vl_logic;
        lsc_prog_incr_cne_cqual: in     vl_logic;
        lsc_prog_incr_cmp_cqual: in     vl_logic;
        nj_cmd_read_com : in     vl_logic;
        nj_cmd_read_dsr : in     vl_logic;
        nj_cmd_prog_com : in     vl_logic;
        j_ins_prog_com  : in     vl_logic;
        jburst_inp      : in     vl_logic;
        dryrun_inp      : in     vl_logic;
        cfg_reset_crc16 : in     vl_logic;
        nj_check_crc    : in     vl_logic;
        decom_last_mask : in     vl_logic;
        dum_dat         : in     vl_logic_vector(7 downto 0);
        jbuf8_rdy       : in     vl_logic;
        jbuf8_dat       : in     vl_logic_vector(7 downto 0);
        njcom_out       : in     vl_logic_vector(7 downto 0);
        dsr_out         : in     vl_logic_vector(7 downto 0);
        wfifo_full      : in     vl_logic;
        rfifo_empty     : in     vl_logic;
        rfifo_out       : in     vl_logic_vector(7 downto 0);
        comp_dic        : in     vl_logic_vector(127 downto 0);
        lsc_sdm         : in     vl_logic;
        dnld_dat        : in     vl_logic_vector(7 downto 0);
        dnld_dat_en     : in     vl_logic;
        lsc_sdm_cfg0    : in     vl_logic;
        lsc_sdm_cfg1    : in     vl_logic;
        sd_authdone_cfg0: in     vl_logic;
        sd_authdone_cfg1: in     vl_logic;
        key_byte        : in     vl_logic_vector(7 downto 0);
        sd_aes_key      : in     vl_logic_vector(255 downto 0);
        sd_auth_en      : in     vl_logic_vector(1 downto 0);
        sd_rand_noise   : in     vl_logic;
        trim_enc_disable: in     vl_logic;
        sd_rand_aes     : in     vl_logic;
        hse_busy        : in     vl_logic_vector(1 downto 0);
        hse_buffer_ready: in     vl_logic;
        hse_pass_fail   : in     vl_logic;
        hse_pf_valid    : in     vl_logic;
        nj_hmac_key     : in     vl_logic;
        nj_hmac_sig     : in     vl_logic;
        nj_ecdsa_key    : in     vl_logic;
        nj_ecdsa_sig    : in     vl_logic;
        njbse_rst_flag  : in     vl_logic;
        lsc_auth_ctrl_cqual: in     vl_logic;
        nj_shf_done     : in     vl_logic;
        nj_last_byte    : in     vl_logic;
        isc_prog_done_c : in     vl_logic;
        njcmd_inf3      : in     vl_logic;
        finish_cdm      : in     vl_logic;
        isc_operational : in     vl_logic;
        ctrl_tran_hse   : in     vl_logic;
        njenable_tran   : in     vl_logic;
        jenable_tran    : in     vl_logic;
        lsc_reset_crc_cq: in     vl_logic;
        bse_sdm_cfg0    : in     vl_logic;
        bse_sdm_cfg1    : in     vl_logic;
        lsc_done_hse    : in     vl_logic;
        njbse_init      : in     vl_logic;
        lsc_reboot_cq   : in     vl_logic;
        sd_uds_trn      : in     vl_logic_vector(127 downto 0);
        uidcode         : in     vl_logic_vector(63 downto 0);
        cdm_done_por    : in     vl_logic;
        hse_trn_out     : in     vl_logic_vector(255 downto 0)
    );
end datap_unit;
