library verilog;
use verilog.vl_types.all;
entity or2x4v1mce is
    port(
        A               : in     vl_logic;
        B               : in     vl_logic;
        Z               : out    vl_logic
    );
end or2x4v1mce;
