library verilog;
use verilog.vl_types.all;
entity cfg_refresh is
    generic(
        INTN_DLY_W      : integer := 4;
        st_idle         : integer := 0;
        st_ppt          : integer := 1;
        st_cdm          : integer := 3;
        st_boot0        : integer := 2;
        st_boot1        : integer := 7;
        st_init         : integer := 5;
        st_boot2        : integer := 4;
        st_exit_accessed: integer := 6
    );
    port(
        ref_ppt         : out    vl_logic;
        ref_cdm         : out    vl_logic;
        ref_init        : out    vl_logic;
        ref_boot0       : out    vl_logic;
        ref_boot1       : out    vl_logic;
        ref_boot2       : out    vl_logic;
        ref_exit        : out    vl_logic;
        initn_tmr       : out    vl_logic;
        exit_accessed   : out    vl_logic;
        ref_sys_slow    : out    vl_logic;
        ref_launch      : out    vl_logic;
        fl_start_ppt    : out    vl_logic;
        fl_start_cdm    : out    vl_logic;
        fl_start_sdm0   : out    vl_logic;
        fl_start_sdm1   : out    vl_logic;
        fl_start_sdm2   : out    vl_logic;
        start_bke       : out    vl_logic;
        ebr_init_en     : out    vl_logic;
        start_bse0      : out    vl_logic;
        start_bse1      : out    vl_logic;
        start_bse2      : out    vl_logic;
        int_prm_nrdy    : out    vl_logic;
        start_wakeup    : out    vl_logic;
        ref_dones       : out    vl_logic_vector(6 downto 0);
        ref_states      : out    vl_logic_vector(6 downto 0);
        wkup_done       : out    vl_logic;
        wkup_done_rise  : out    vl_logic;
        rst_wkup_done   : out    vl_logic;
        rst_ctrl01_onfail: out    vl_logic;
        fl_start_sdm_cfg0: out    vl_logic;
        fl_start_sdm_cfg1: out    vl_logic;
        wkup_to_reboot  : out    vl_logic;
        wkup_to_reboot_st: out    vl_logic;
        cdm_done_por    : out    vl_logic;
        HFC_EN          : in     vl_logic;
        hfc_select_pin  : in     vl_logic;
        scanen          : in     vl_logic;
        smclk           : in     vl_logic;
        por             : in     vl_logic;
        fsafe           : in     vl_logic;
        ref_rst_sync    : in     vl_logic;
        isc_nj_enabled  : in     vl_logic;
        exit_fl_offline_exec: in     vl_logic;
        exit_normal_exec: in     vl_logic;
        fsd_persist_initn: in     vl_logic;
        programn_pin_sync: in     vl_logic;
        initn_pin_sync  : in     vl_logic;
        p_eboot0p       : in     vl_logic;
        p_eboot1p       : in     vl_logic;
        p_eboot1s       : in     vl_logic;
        p_eboot2p       : in     vl_logic;
        p_eboot2s       : in     vl_logic;
        p_nboot         : in     vl_logic;
        p_iboot0p       : in     vl_logic;
        p_iboot1p       : in     vl_logic;
        p_iboot1s       : in     vl_logic;
        p_iboot2p       : in     vl_logic;
        p_iboot2s       : in     vl_logic;
        ctrl_ncdm       : in     vl_logic;
        ctrl_nbke       : in     vl_logic;
        ctrl_ebr_init_en: in     vl_logic;
        ctrl_hfc_hd     : in     vl_logic;
        isc_done        : in     vl_logic;
        access_sram     : in     vl_logic;
        access_flash    : in     vl_logic;
        enter_offline_exec: in     vl_logic;
        enter_offline_eqv: in     vl_logic;
        ref_start       : in     vl_logic;
        jaccessed_sync  : in     vl_logic;
        finish_ppt      : in     vl_logic;
        finish_cdm      : in     vl_logic;
        finish_sdm      : in     vl_logic;
        finish_bke      : in     vl_logic;
        finish_bse      : in     vl_logic;
        njbse_finish    : in     vl_logic;
        fail_sdm_a      : in     vl_logic;
        fail_sdm_b      : in     vl_logic;
        fail_bse        : in     vl_logic;
        wkup_done_cib   : in     vl_logic;
        flash_done_a    : in     vl_logic;
        flash_done_b    : in     vl_logic;
        p_iboot0s       : in     vl_logic;
        finish_auth     : in     vl_logic;
        fail_auth       : in     vl_logic;
        reset_auth      : in     vl_logic;
        auth_en         : in     vl_logic;
        auth_ready      : in     vl_logic;
        dec_ready       : in     vl_logic;
        tc_to_reboot_en : in     vl_logic;
        tc_to           : in     vl_logic;
        tc_to_reboot_mode: in     vl_logic;
        bse_timeout_err : in     vl_logic;
        vrbp_auth_done  : in     vl_logic
    );
end cfg_refresh;
