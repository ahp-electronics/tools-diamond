--
@ER--B$FbsEHo0OR52gR4g-cRRj.jd$R1MHbDO$H0ROQM
R--fN]C8:CsR#//$DMbH0OH$N/lb..jjDjdNl0/NCbbsN#/0D0/HoL/CFM_s.ONNN/slI_s38PEyf4R

--
-
-
R--1bHlD)CRqIvRHR0E#oHMDqCR7 7)1V1RFLsRFR0Es8CNR8NMRHIs0-C
-NRas0oCRp:RkMOC0RR-mq)BR
.q---
-D

HNLssH$RC;CC
Ck#RCHCC03#8F_Do_HO4c4n3DND;#
kCCRHC#C30D8_FOoH_o#HM3C8N;DD
LDHs$NsROFsN
.;kR#CFNsO.s3FOFNOlNb3D
D;CHM00)$Rq)v_W#RH
RRRRMoCCOsHRR5
RRRRRVRRNDlH$#:R0MsHo=R:RF"MM;C"
RRRRRRRR8IH0:ERR0HMCsoCRR:=4
;RRRRRRRRRNs88I0H8ERR:HCM0oRCs:c=R;RRRRRRRRR--LRHoCkMFoVERF8sRCEb0
RRRRRRRRb8C0:ERR0HMCsoCRR:=R;4n
RRRRRRRRk8F0C_soRR:LDFFCRNM:V=RNCD#;RRRR-R-R#ENR0FkbRk0s
CoRRRRRRRR8_HMsRCo:FRLFNDCM=R:RDVN#RC;RRRRRR--ERN#8NN0RbHMks0RCRo
RRRRRNRR8_8ssRCo:FRLFNDCM=R:RDVN#RCRRRRR-E-RNN8R8C8s#s#RCRo
RRRRR2RR;R
RRFRbs50R
RRRRRRRRz7maRR:FRk0#_08DHFoOC_POs0F58IH04E-RI8FMR0Fj
2;RRRRRRRR7RQhRH:RM0R#8F_Do_HOP0COFIs5HE80-84RF0IMF2Rj;R
RRRRRR7Rq7:)RRRHM#_08DHFoOC_POs0F58N8s8IH04E-RI8FMR0Fj
2;RRRRRRRRWR R:MRHR8#0_oDFHRO;RRRRR-R-RHIs0CCRMDNLCFRVsNRslR
RRRRRRpRBiRR:H#MR0D8_FOoH;RRRRRRR-O-RD	FORsVFRlsN,8RN8Rs,8
HMRRRRRRRRmiBpRH:RM0R#8F_DoRHORRRRR-R-R0FbRFODOV	RF8sRF
k0RRRRRRRR2C;
MC8RM00H$qR)vW_);-

--
-RswH#H0RlCbDl0CMNF0HMkRl#L0RCNROD8DCRONsE-j
-s
NO0EHCkO0sNCRsjOERRFV)_qv)HWR#F
OMN#0MM0RkOl_C#DD_C8CbRR:HCM0oRCs:5=R5b8C0-ERR/424;n2RRRRR-RR-RRyFsVRFRI#F)VRBnw4XRcZODCD#CRMC88C
MOF#M0N0kRMlC_OD_D#ICH8RH:RMo0CC:sR=5R5I0H8ERR-4c2/2R;RRRRRR-R-RFyRVFRODMkl#VRFRw)B4cnXZCRODRD#M8CCC-8
-b0$CkRF0k_L#$_0bHCR#sRNsRN$5lMk_DOCD8#RF0IMF,RjR8IH04E-RI8FMR0FjF2RV0R#8F_Do;HO
#--HNoMDkRF0k_L#RR:F_k0L_k#0C$b;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-.-R7sRNsRN$F8VRFRk05bHMk00RFsR0H0-#N#0C2H
#oDMNR0Fk_RCM:0R#8F_Do_HOP0COFMs5kOl_C#DD_C8CbFR8IFM0R;j2RRRRRRRR-C-RMDNLCV#RF0sRs#H-0CN0#H
#oDMNRCIb_RCM:0R#8F_Do_HOP0COFMs5kOl_C#DD_C8CbFR8IFM0R;j2RRRRRRRR-I-RsCH0RNCML#DCRsVFROCNEFRsIVRFRv)qRDOCD##
HNoMDMRH_osCR#:R0D8_FOoH_OPC05FsI0H8ER+d8MFI0jFR2R;RRRRRRRRR-k-R#RC80sFRC#oH0RCs7RQh
o#HMRNDF_k0sRCo:0R#8F_Do_HOP0COFIs5HE80+8dRF0IMF2Rj;RRRRRRRR-R-RCk#8FR0RosCHC#0smR7z#a
HNoMD8RN_osCR#:R0D8_FOoH_OPC05FsNs88I0H8ER-48MFI0jFR2R;RRRRR-k-R#RC80sFRC#oH0RCsq)77
o#HMRNDD_FINs88R#:R0D8_FOoH_OPC05FsdFR8IFM0R;j2RRRRRRRRRRRRR-R-R8N8sHRL0H#RM0bkRR0F)RqvODCD#cR5R0LH#CRsJskHC
82
oLCH
M
RRRR-Q-RV8RN8HsI8R0E<RRcNH##o'MRj0'RFMRkk8#CR0LH#R
RR4RzRRR:H5VRNs88I0H8ERR=4o2RCsMCN
0CRRRRRRRRD_FINs88RR<="jjj"RR&Ns8_Cjo52R;
RCRRMo8RCsMCNR0Cz
4;RRRRzR.R:VRHR85N8HsI8R0E=2R.RMoCC0sNCR
RRRRRRFRDI8_N8<sR=jR"j&"RR_N8s5Co4FR8IFM0R;j2
RRRR8CMRMoCC0sNC.Rz;R
RRdRzRRR:H5VRNs88I0H8ERR=do2RCsMCN
0CRRRRRRRRD_FINs88RR<='Rj'&8RN_osC58.RF0IMF2Rj;R
RRMRC8CRoMNCs0zCRdR;
RzRRc:RRRRHV58N8s8IH0>ERRRd2oCCMsCN0
RRRRRRRRIDF_8N8s=R<R_N8s5CodFR8IFM0R;j2
RRRR8CMRMoCC0sNCcRz;R

R-RR-VRQRH58MC_sos2RC#oH0RCs7RQhkM#HopRBiR
RR6RzRRR:H5VR8_HMs2CoRMoCC0sNCR
RRRRRRsRbF#OC#BR5pRi,72QhRoLCHRM
RRRRRRRRRHRRVBR5p=iRR''4R8NMRiBp'CCPMR020MEC
RRRRRRRRRRRRRRRR_HMsRCo<5=R"jjjj&"RRh7Q2R;
RRRRRRRRRCRRMH8RVR;
RRRRRCRRMb8RsCFO#
#;RRRRCRM8oCCMsCN0R;z6
RRRRRznRH:RVMR5F80RHsM_CRo2oCCMsCN0
RRRRRRRRRRRR_HMsRCo<5=R"jjjj&"RRh7Q2R;
RCRRMo8RCsMCNR0Cz
n;
RRRRR--Q5VR80Fk_osC2CRso0H#C7sRmRzakM#HoBRmpRi
RzRR(:RRRRHV5k8F0C_soo2RCsMCN
0CRRRRRRRRbOsFCR##5pmBiF,Rks0_CRo2LHCoMR
RRRRRRRRRRVRHRB5mp=iRR''4R8NMRpmBiP'CC2M0RC0EMR
RRRRRRRRRRRRRRmR7z<aR=kRF0C_soH5I8-0E4FR8IFM0R;j2
RRRRRRRRRRRR8CMR;HV
RRRRRRRR8CMRFbsO#C#;R
RRRRRRMRC8CRoMNCs0zCR(R;
RzRRU:RRRRHV50MFRk8F0C_soo2RCsMCN
0CRRRRRRRRRRRR7amzRR<=F_k0s5CoI0H8ER-48MFI0jFR2R;
RCRRMo8RCsMCNR0Cz
U;
RRRRR--Q5VRNs88_osC2CRso0H#CqsR7R7)kM#HopRBiR
RRgRzRRR:H5VRNs88_osC2CRoMNCs0RC
RRRRRbRRsCFO#5#RB,piR7q7)L2RCMoH
RRRRRRRRRRRRRHV5iBpR'=R4N'RMB8RpCi'P0CM2ER0CRM
RRRRRRRRRRRRRNRR8C_so=R<R7q7)85N8HsI8-0E4FR8IFM0R;j2
RRRRRRRRRRRR8CMR;HV
RRRRRRRR8CMRFbsO#C#;R
RRMRC8CRoMNCs0zCRgR;
RzRR4:jRRRHV50MFR8N8sC_soo2RCsMCN
0CRRRRRRRRRRRRNs8_C<oR=7Rq7
);RRRRCRM8oCCMsCN0Rjz4;R
RRRRRRRR
R-RR-CRtMNCs00CRE)CRqOvRC#DDR8NMRD#CCRO0DHFoOR
RR4Rz4RR:VRFsHMRHRlMk_DOCD8#_CRCb8MFI0jFRRMoCC0sNCR
RR-R-RRQV58N8s8IH0>ERRRc2M8CCRR0FONsC0ICRsCH0RNCMLRDCNRM8Fbk0kC0RMDNLCCR#D0CORoDFHRO
RRRRRzRR4:.RRRHV58N8s8IH0>ERRRc2oCCMsCN0
RRRRRRRRRRRRRRRR0Fk_5CMH<2R=jR''ERIC5MRNs8_CNo58I8sHE80-84RF0IMF2RcRH=R2DRC#'CR4
';RRRRRRRRRRRRRRRRI_bCCHM52=R<R''4RCIEMNR58C_so85N8HsI8-0E4FR8IFM0RRc2=2RHR#CDCjR''R;
RRRRRRRRRCRRMo8RCsMCNR0Cz;4.
RRRRR--Q5VRNs88I0H8E=R<RRc2MIFRsCH0RNCMLRDCFFsRkk0b0MRCNCLDRD#CCRO0DHFoOCRMC88C
RRRRdz4RH:RVNR58I8sHE80RR<=co2RCsMCN
0CRRRRRRRRRRRRF_k0CHM52=R<R''j;R
RRRRRRRRRRRRRRbRICM_C5RH2<'=R4
';RRRRRRRRRRRRCRM8oCCMsCN0Rdz4;R
RR-R-RCtMsCN0RC0ERv)qRDOCDI#RHR0E0-sH#00NCR#
RRRRRzRR4:cRRsVFRH[RMkRMlC_OD_D#ICH8RI8FMR0FjCRoMNCs0RC
RRRRRRRRRzRR):qvRw)B4cnXZRR
RRRRRRRRRbRRFRs0lRNb5Qa)RR=>F_k0CHM527,RQ=jR>MRH_osC5*5c[,22R47QRR=>HsM_C5o5c2*[+,42R.7QRR=>HsM_C5o5c2*[+,.2RR
RRRRRRRRRRRRRRRRRRRRRRRRR7RQd=H>RMC_soc55*+[2dR2,qR7j=D>RFNI_858sjR2,qR74=D>RFNI_858s4R2,qR7.=D>RFNI_858s.
2,RRRRRRRRRRRRRRRRRRRRRRRRR7Rqd>R=RIDF_8N8s25d,)RW =hR> RW,uRW >R=RCIb_5CMHR2,B=iR>pRBi7,Rm=jR>kRF0C_so[55*2c2,R
RRRRRRRRRRRRRRRRRRRRRRRRR7Rm4=F>Rks0_C5o5[2*c+,42R.7mRR=>F_k0s5Co5c[*22+.,mR7d>R=R0Fk_osC5*5[cd2+2
2;RRRRRRRRRRRRCRM8oCCMsCN0Rcz4;R
RRRRRRMRC8CRoMNCs0zCR4
4;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRM
C8sRNO0EHCkO0sNCRsjOE;



