library verilog;
use verilog.vl_types.all;
entity fx65_osc_1inv is
    port(
        \in\            : in     vl_logic;
        \out\           : out    vl_logic
    );
end fx65_osc_1inv;
