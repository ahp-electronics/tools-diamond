library verilog;
use verilog.vl_types.all;
entity cfg is
    generic(
        MASTER_SERI     : integer := 8;
        MASTER_PARA     : integer := 12;
        ASYNC_PERI      : integer := 13;
        SLAVE_SERI      : integer := 15;
        SLAVE_PARA      : integer := 9;
        FPSC_PARA       : integer := 7;
        MASTER_BYTE     : integer := 6;
        FLASH_SPI03     : integer := 5;
        FLASH_SPIX      : integer := 4;
        MPC_BYTE        : integer := 10;
        MPC_HWORD       : integer := 11;
        MPC_WORD        : integer := 14;
        CHK_PRE         : integer := 0;
        CHK_ID          : integer := 1;
        CHK_HDR         : integer := 2;
        CHK_FPGA        : integer := 3;
        CHK_RAM         : integer := 6;
        CHK_FPSC        : integer := 5;
        CHK_POST        : integer := 7
    );
    port(
        CODE0           : in     vl_logic_vector(7 downto 0);
        CODE1           : in     vl_logic_vector(7 downto 0);
        CODE2           : in     vl_logic_vector(7 downto 0);
        CODE3           : in     vl_logic_vector(7 downto 0);
        CODE4           : in     vl_logic_vector(7 downto 0);
        CODE5           : in     vl_logic_vector(7 downto 0);
        CODE6           : in     vl_logic_vector(7 downto 0);
        CODE7           : in     vl_logic_vector(7 downto 0);
        EN_COUNT6       : in     vl_logic;
        LAST_ADDR       : in     vl_logic_vector(13 downto 0);
        PARTID          : in     vl_logic_vector(31 downto 12);
        HGRANT_CFG      : in     vl_logic;
        HREADY_CFG      : in     vl_logic;
        HRESET_N        : in     vl_logic;
        HRESP_CFG       : in     vl_logic_vector(1 downto 0);
        REPEAT_RDBK     : in     vl_logic;
        MPI_USR_ENABLE  : in     vl_logic;
        SYS_RD_CFG      : in     vl_logic;
        SYS_GSR         : in     vl_logic;
        PRGM_MPI        : in     vl_logic;
        PRGM_FPSC       : in     vl_logic;
        PRGM_USER       : in     vl_logic;
        SYS_DAISY       : in     vl_logic;
        RDATA_ACK       : in     vl_logic;
        WDATA_READY     : in     vl_logic;
        RDATA_SIZE      : in     vl_logic_vector(1 downto 0);
        WDATA_SIZE      : in     vl_logic_vector(1 downto 0);
        WDATA           : in     vl_logic_vector(31 downto 0);
        RDBK_ADDR       : in     vl_logic_vector(13 downto 0);
        MPI_RD_DATA     : in     vl_logic_vector(7 downto 3);
        MPI_TRI_DATA    : in     vl_logic;
        MPI_TRI_CNTL    : in     vl_logic;
        RCLKS           : in     vl_logic;
        HCLK            : in     vl_logic;
        CCLK            : in     vl_logic;
        SER_CCLK        : in     vl_logic;
        CFG_CK          : in     vl_logic;
        OSC_DIV128      : in     vl_logic;
        J_SPI_PROG      : in     vl_logic;
        J_SHDR          : in     vl_logic;
        J_SCANIN        : in     vl_logic;
        J_TCK           : in     vl_logic;
        PRGM_JTAG       : in     vl_logic;
        RD_CFG_JTAG     : in     vl_logic;
        TDI_JTAG        : in     vl_logic;
        BS_MODE         : in     vl_logic;
        SCAN_CFG        : in     vl_logic;
        CFG_PRGM_N      : in     vl_logic;
        CFG_RESET_N     : in     vl_logic;
        RD_CFG          : in     vl_logic;
        PWRUP_E9        : in     vl_logic;
        PWRUP_NPUR      : in     vl_logic;
        ADDR_HIGH_DEL_N : in     vl_logic;
        RDBK_ZERO_ALL_N : in     vl_logic;
        DEL_D           : in     vl_logic_vector(7 downto 0);
        RDBK_DOUT       : in     vl_logic_vector(7 downto 0);
        PTEST_N         : in     vl_logic;
        DONEIN          : in     vl_logic;
        INITIN_N        : in     vl_logic;
        CS0_N           : in     vl_logic;
        CS1             : in     vl_logic;
        RD_N            : in     vl_logic;
        WR_N            : in     vl_logic;
        MODE            : in     vl_logic_vector(3 downto 0);
        SPI_ADDR_RAM    : in     vl_logic_vector(31 downto 0);
        EN_SPI_RAM_N    : in     vl_logic;
        EN_SED_RAM      : in     vl_logic;
        RDBK_REG_RAM    : in     vl_logic;
        MPI_RST_RAM     : in     vl_logic;
        SYS_RST_RAM     : in     vl_logic;
        MPI_ASYNC_RAM   : in     vl_logic;
        GSRN_SYNC_RAM   : in     vl_logic;
        RST_GSRN_RAM    : in     vl_logic;
        GSRN_INV_RAM    : in     vl_logic;
        OSC_DIV_RAM     : in     vl_logic_vector(2 downto 0);
        MPI_CLK_RAM     : in     vl_logic;
        FPSC_CLK_RAM    : in     vl_logic;
        USR_CLK_RAM     : in     vl_logic;
        OSC_CLK_RAM     : in     vl_logic;
        DIS_MODES_RAM   : in     vl_logic;
        EN_OSC_RAM      : in     vl_logic;
        EXT_CCLK_RAM    : in     vl_logic;
        TEST_CTR_RAM    : in     vl_logic;
        RST_BUS_RAM_N   : in     vl_logic;
        RST_HCLK_RAM_N  : in     vl_logic;
        RST_RAM_RAM_N   : in     vl_logic;
        SCLK_RAM        : in     vl_logic;
        EN_CAPTURE_RAM  : in     vl_logic;
        EN_ONCE_RAM     : in     vl_logic;
        EN_RDBK_RAM     : in     vl_logic;
        EN_READCAP_RAM  : in     vl_logic;
        EN_MPI_PARITY_RAM: in     vl_logic;
        MODE_RAM        : in     vl_logic_vector(3 downto 0);
        DONE_RAM        : in     vl_logic_vector(1 downto 0);
        STRT_RAM        : in     vl_logic_vector(4 downto 0);
        TRI_RAM         : in     vl_logic_vector(3 downto 0);
        RD_CFG_USR      : in     vl_logic;
        MPI_RST_N       : in     vl_logic;
        SYS_RST_N       : in     vl_logic;
        USR_START_CLK   : in     vl_logic;
        USR_GSR         : in     vl_logic;
        CAPT_I_N        : in     vl_logic;
        FPSC_GSR        : in     vl_logic;
        HBUSREQ_CFG     : out    vl_logic;
        HLOCK_CFG       : out    vl_logic;
        HWRITE_CFG      : out    vl_logic;
        HBURST_CFG      : out    vl_logic;
        HTRANS_CFG      : out    vl_logic_vector(1 downto 0);
        HSIZE_CFG       : out    vl_logic_vector(1 downto 0);
        HADDR_CFG       : out    vl_logic_vector(17 downto 0);
        HWDATA_CFG      : out    vl_logic_vector(35 downto 0);
        RFR_SEL         : out    vl_logic_vector(3 downto 0);
        HRESET_OUT      : out    vl_logic;
        HCLK_SWITCH     : out    vl_logic;
        RST_LOCK        : out    vl_logic;
        RDATA_READY     : out    vl_logic;
        WDATA_ACK       : out    vl_logic;
        CFG_IRQ_DATA    : out    vl_logic;
        FPSC_BIT_ERR    : out    vl_logic;
        RAM_BIT_ERR     : out    vl_logic;
        RDBK_ADDR_ERR   : out    vl_logic;
        BUS_DATA_LOST   : out    vl_logic;
        BUS_TRAP_ADDR   : out    vl_logic_vector(17 downto 0);
        CFG_BUS_ERR     : out    vl_logic_vector(1 downto 0);
        BUS_ERR_ADDR    : out    vl_logic_vector(17 downto 0);
        ERR_FLAG        : out    vl_logic_vector(1 downto 0);
        RDATA           : out    vl_logic_vector(31 downto 0);
        MPI_DATA_PORT   : out    vl_logic_vector(2 downto 0);
        MPI_DP_ENABLE   : out    vl_logic;
        MPI_SYNC        : out    vl_logic;
        MPI_RESET_N     : out    vl_logic;
        OSC_DIV_EN      : out    vl_logic;
        HCLK_SEL        : out    vl_logic_vector(2 downto 0);
        SCLK_SEL        : out    vl_logic_vector(1 downto 0);
        CCLK_SEL        : out    vl_logic_vector(1 downto 0);
        CK_SEL          : out    vl_logic_vector(2 downto 0);
        CFGDOUT_JTAG_N  : out    vl_logic;
        BS_RST_JTAG_N   : out    vl_logic;
        EN_OSC          : out    vl_logic;
        PWR_ON          : out    vl_logic;
        EN_ADDR         : out    vl_logic;
        RST_ADDR_REG    : out    vl_logic;
        GOT_ADDR        : out    vl_logic;
        EN_ADDR_INCR    : out    vl_logic;
        SHIFT_ADDR_1ST  : out    vl_logic;
        SHIFT_ADDR_2ND  : out    vl_logic;
        RST_DATA_REG_N  : out    vl_logic;
        GOT_DATA        : out    vl_logic;
        INIT_1_DATA     : out    vl_logic;
        CFG_DATA_WR     : out    vl_logic;
        SERIAL_DATA     : out    vl_logic;
        LD_RDBKD        : out    vl_logic;
        CFG_DATA_PC     : out    vl_logic;
        CFG_DATA        : out    vl_logic_vector(7 downto 0);
        PAD_DONE        : out    vl_logic;
        INIT_N          : out    vl_logic;
        HDC             : out    vl_logic;
        LDC_N           : out    vl_logic;
        RDY_BUSY_N      : out    vl_logic;
        DOUT            : out    vl_logic;
        QOUT            : out    vl_logic;
        RDBK_DATA       : out    vl_logic;
        RDBK_TDO_EN     : out    vl_logic;
        PD_OUT          : out    vl_logic_vector(7 downto 3);
        PA_OUT          : out    vl_logic_vector(21 downto 0);
        EN_CCLK_N       : out    vl_logic;
        PD7_3_TS        : out    vl_logic;
        PRDY_TS         : out    vl_logic;
        PD2_0_TS        : out    vl_logic;
        PD15_8_TS       : out    vl_logic;
        PD31_16_TS      : out    vl_logic;
        MPI_CNTL_TS     : out    vl_logic;
        MPI_DP_TS       : out    vl_logic_vector(2 downto 0);
        MPI_DP_TRI_ION  : out    vl_logic_vector(2 downto 0);
        MPI_TRI_ION     : out    vl_logic_vector(2 downto 0);
        ADDR_TS         : out    vl_logic;
        SPI_TRI_ION     : out    vl_logic;
        DEBUG_BUS       : out    vl_logic_vector(15 downto 0);
        CAPTURE         : out    vl_logic;
        TRI_ION         : out    vl_logic;
        DONE            : out    vl_logic;
        GSR_N           : out    vl_logic;
        GSRN_SYNC       : out    vl_logic;
        EN_PDWN         : out    vl_logic;
        PWRUPRES        : out    vl_logic;
        PAD_INIT_N      : out    vl_logic
    );
end cfg;
