library verilog;
use verilog.vl_types.all;
entity PCSD_sim is
    generic(
        CONFIG_FILE     : string  := "configfile.txt";
        QUAD_MODE       : string  := "SINGLE";
        PLL_SRC         : string  := "REFCLK_EXT";
        CH0_CDR_SRC     : string  := "REFCLK_EXT";
        CH1_CDR_SRC     : string  := "REFCLK_EXT";
        CH2_CDR_SRC     : string  := "REFCLK_EXT";
        CH3_CDR_SRC     : string  := "REFCLK_EXT"
    );
    port(
        HDINN0          : in     vl_logic;
        HDINN1          : in     vl_logic;
        HDINN2          : in     vl_logic;
        HDINN3          : in     vl_logic;
        HDINP0          : in     vl_logic;
        HDINP1          : in     vl_logic;
        HDINP2          : in     vl_logic;
        HDINP3          : in     vl_logic;
        REFCLKN         : in     vl_logic;
        REFCLKP         : in     vl_logic;
        CIN0            : in     vl_logic;
        CIN1            : in     vl_logic;
        CIN2            : in     vl_logic;
        CIN3            : in     vl_logic;
        CIN4            : in     vl_logic;
        CIN5            : in     vl_logic;
        CIN6            : in     vl_logic;
        CIN7            : in     vl_logic;
        CIN8            : in     vl_logic;
        CIN9            : in     vl_logic;
        CIN10           : in     vl_logic;
        CIN11           : in     vl_logic;
        CYAWSTN         : in     vl_logic;
        FF_EBRD_CLK_0   : in     vl_logic;
        FF_EBRD_CLK_1   : in     vl_logic;
        FF_EBRD_CLK_2   : in     vl_logic;
        FF_EBRD_CLK_3   : in     vl_logic;
        FF_RXI_CLK_0    : in     vl_logic;
        FF_RXI_CLK_1    : in     vl_logic;
        FF_RXI_CLK_2    : in     vl_logic;
        FF_RXI_CLK_3    : in     vl_logic;
        FF_TX_D_0_0     : in     vl_logic;
        FF_TX_D_0_1     : in     vl_logic;
        FF_TX_D_0_2     : in     vl_logic;
        FF_TX_D_0_3     : in     vl_logic;
        FF_TX_D_0_4     : in     vl_logic;
        FF_TX_D_0_5     : in     vl_logic;
        FF_TX_D_0_6     : in     vl_logic;
        FF_TX_D_0_7     : in     vl_logic;
        FF_TX_D_0_8     : in     vl_logic;
        FF_TX_D_0_9     : in     vl_logic;
        FF_TX_D_0_10    : in     vl_logic;
        FF_TX_D_0_11    : in     vl_logic;
        FF_TX_D_0_12    : in     vl_logic;
        FF_TX_D_0_13    : in     vl_logic;
        FF_TX_D_0_14    : in     vl_logic;
        FF_TX_D_0_15    : in     vl_logic;
        FF_TX_D_0_16    : in     vl_logic;
        FF_TX_D_0_17    : in     vl_logic;
        FF_TX_D_0_18    : in     vl_logic;
        FF_TX_D_0_19    : in     vl_logic;
        FF_TX_D_0_20    : in     vl_logic;
        FF_TX_D_0_21    : in     vl_logic;
        FF_TX_D_0_22    : in     vl_logic;
        FF_TX_D_0_23    : in     vl_logic;
        FF_TX_D_1_0     : in     vl_logic;
        FF_TX_D_1_1     : in     vl_logic;
        FF_TX_D_1_2     : in     vl_logic;
        FF_TX_D_1_3     : in     vl_logic;
        FF_TX_D_1_4     : in     vl_logic;
        FF_TX_D_1_5     : in     vl_logic;
        FF_TX_D_1_6     : in     vl_logic;
        FF_TX_D_1_7     : in     vl_logic;
        FF_TX_D_1_8     : in     vl_logic;
        FF_TX_D_1_9     : in     vl_logic;
        FF_TX_D_1_10    : in     vl_logic;
        FF_TX_D_1_11    : in     vl_logic;
        FF_TX_D_1_12    : in     vl_logic;
        FF_TX_D_1_13    : in     vl_logic;
        FF_TX_D_1_14    : in     vl_logic;
        FF_TX_D_1_15    : in     vl_logic;
        FF_TX_D_1_16    : in     vl_logic;
        FF_TX_D_1_17    : in     vl_logic;
        FF_TX_D_1_18    : in     vl_logic;
        FF_TX_D_1_19    : in     vl_logic;
        FF_TX_D_1_20    : in     vl_logic;
        FF_TX_D_1_21    : in     vl_logic;
        FF_TX_D_1_22    : in     vl_logic;
        FF_TX_D_1_23    : in     vl_logic;
        FF_TX_D_2_0     : in     vl_logic;
        FF_TX_D_2_1     : in     vl_logic;
        FF_TX_D_2_2     : in     vl_logic;
        FF_TX_D_2_3     : in     vl_logic;
        FF_TX_D_2_4     : in     vl_logic;
        FF_TX_D_2_5     : in     vl_logic;
        FF_TX_D_2_6     : in     vl_logic;
        FF_TX_D_2_7     : in     vl_logic;
        FF_TX_D_2_8     : in     vl_logic;
        FF_TX_D_2_9     : in     vl_logic;
        FF_TX_D_2_10    : in     vl_logic;
        FF_TX_D_2_11    : in     vl_logic;
        FF_TX_D_2_12    : in     vl_logic;
        FF_TX_D_2_13    : in     vl_logic;
        FF_TX_D_2_14    : in     vl_logic;
        FF_TX_D_2_15    : in     vl_logic;
        FF_TX_D_2_16    : in     vl_logic;
        FF_TX_D_2_17    : in     vl_logic;
        FF_TX_D_2_18    : in     vl_logic;
        FF_TX_D_2_19    : in     vl_logic;
        FF_TX_D_2_20    : in     vl_logic;
        FF_TX_D_2_21    : in     vl_logic;
        FF_TX_D_2_22    : in     vl_logic;
        FF_TX_D_2_23    : in     vl_logic;
        FF_TX_D_3_0     : in     vl_logic;
        FF_TX_D_3_1     : in     vl_logic;
        FF_TX_D_3_2     : in     vl_logic;
        FF_TX_D_3_3     : in     vl_logic;
        FF_TX_D_3_4     : in     vl_logic;
        FF_TX_D_3_5     : in     vl_logic;
        FF_TX_D_3_6     : in     vl_logic;
        FF_TX_D_3_7     : in     vl_logic;
        FF_TX_D_3_8     : in     vl_logic;
        FF_TX_D_3_9     : in     vl_logic;
        FF_TX_D_3_10    : in     vl_logic;
        FF_TX_D_3_11    : in     vl_logic;
        FF_TX_D_3_12    : in     vl_logic;
        FF_TX_D_3_13    : in     vl_logic;
        FF_TX_D_3_14    : in     vl_logic;
        FF_TX_D_3_15    : in     vl_logic;
        FF_TX_D_3_16    : in     vl_logic;
        FF_TX_D_3_17    : in     vl_logic;
        FF_TX_D_3_18    : in     vl_logic;
        FF_TX_D_3_19    : in     vl_logic;
        FF_TX_D_3_20    : in     vl_logic;
        FF_TX_D_3_21    : in     vl_logic;
        FF_TX_D_3_22    : in     vl_logic;
        FF_TX_D_3_23    : in     vl_logic;
        FF_TXI_CLK_0    : in     vl_logic;
        FF_TXI_CLK_1    : in     vl_logic;
        FF_TXI_CLK_2    : in     vl_logic;
        FF_TXI_CLK_3    : in     vl_logic;
        FFC_CK_CORE_RX_0: in     vl_logic;
        FFC_CK_CORE_RX_1: in     vl_logic;
        FFC_CK_CORE_RX_2: in     vl_logic;
        FFC_CK_CORE_RX_3: in     vl_logic;
        FFC_CK_CORE_TX  : in     vl_logic;
        FFC_EI_EN_0     : in     vl_logic;
        FFC_EI_EN_1     : in     vl_logic;
        FFC_EI_EN_2     : in     vl_logic;
        FFC_EI_EN_3     : in     vl_logic;
        FFC_ENABLE_CGALIGN_0: in     vl_logic;
        FFC_ENABLE_CGALIGN_1: in     vl_logic;
        FFC_ENABLE_CGALIGN_2: in     vl_logic;
        FFC_ENABLE_CGALIGN_3: in     vl_logic;
        FFC_FB_LOOPBACK_0: in     vl_logic;
        FFC_FB_LOOPBACK_1: in     vl_logic;
        FFC_FB_LOOPBACK_2: in     vl_logic;
        FFC_FB_LOOPBACK_3: in     vl_logic;
        FFC_LANE_RX_RST_0: in     vl_logic;
        FFC_LANE_RX_RST_1: in     vl_logic;
        FFC_LANE_RX_RST_2: in     vl_logic;
        FFC_LANE_RX_RST_3: in     vl_logic;
        FFC_LANE_TX_RST_0: in     vl_logic;
        FFC_LANE_TX_RST_1: in     vl_logic;
        FFC_LANE_TX_RST_2: in     vl_logic;
        FFC_LANE_TX_RST_3: in     vl_logic;
        FFC_MACRO_RST   : in     vl_logic;
        FFC_PCI_DET_EN_0: in     vl_logic;
        FFC_PCI_DET_EN_1: in     vl_logic;
        FFC_PCI_DET_EN_2: in     vl_logic;
        FFC_PCI_DET_EN_3: in     vl_logic;
        FFC_PCIE_CT_0   : in     vl_logic;
        FFC_PCIE_CT_1   : in     vl_logic;
        FFC_PCIE_CT_2   : in     vl_logic;
        FFC_PCIE_CT_3   : in     vl_logic;
        FFC_PFIFO_CLR_0 : in     vl_logic;
        FFC_PFIFO_CLR_1 : in     vl_logic;
        FFC_PFIFO_CLR_2 : in     vl_logic;
        FFC_PFIFO_CLR_3 : in     vl_logic;
        FFC_QUAD_RST    : in     vl_logic;
        FFC_RRST_0      : in     vl_logic;
        FFC_RRST_1      : in     vl_logic;
        FFC_RRST_2      : in     vl_logic;
        FFC_RRST_3      : in     vl_logic;
        FFC_RXPWDNB_0   : in     vl_logic;
        FFC_RXPWDNB_1   : in     vl_logic;
        FFC_RXPWDNB_2   : in     vl_logic;
        FFC_RXPWDNB_3   : in     vl_logic;
        FFC_SB_INV_RX_0 : in     vl_logic;
        FFC_SB_INV_RX_1 : in     vl_logic;
        FFC_SB_INV_RX_2 : in     vl_logic;
        FFC_SB_INV_RX_3 : in     vl_logic;
        FFC_SB_PFIFO_LP_0: in     vl_logic;
        FFC_SB_PFIFO_LP_1: in     vl_logic;
        FFC_SB_PFIFO_LP_2: in     vl_logic;
        FFC_SB_PFIFO_LP_3: in     vl_logic;
        FFC_SIGNAL_DETECT_0: in     vl_logic;
        FFC_SIGNAL_DETECT_1: in     vl_logic;
        FFC_SIGNAL_DETECT_2: in     vl_logic;
        FFC_SIGNAL_DETECT_3: in     vl_logic;
        FFC_SYNC_TOGGLE : in     vl_logic;
        FFC_TRST        : in     vl_logic;
        FFC_TXPWDNB_0   : in     vl_logic;
        FFC_TXPWDNB_1   : in     vl_logic;
        FFC_TXPWDNB_2   : in     vl_logic;
        FFC_TXPWDNB_3   : in     vl_logic;
        FFC_RATE_MODE_RX_0: in     vl_logic;
        FFC_RATE_MODE_RX_1: in     vl_logic;
        FFC_RATE_MODE_RX_2: in     vl_logic;
        FFC_RATE_MODE_RX_3: in     vl_logic;
        FFC_RATE_MODE_TX_0: in     vl_logic;
        FFC_RATE_MODE_TX_1: in     vl_logic;
        FFC_RATE_MODE_TX_2: in     vl_logic;
        FFC_RATE_MODE_TX_3: in     vl_logic;
        FFC_DIV11_MODE_RX_0: in     vl_logic;
        FFC_DIV11_MODE_RX_1: in     vl_logic;
        FFC_DIV11_MODE_RX_2: in     vl_logic;
        FFC_DIV11_MODE_RX_3: in     vl_logic;
        FFC_DIV11_MODE_TX_0: in     vl_logic;
        FFC_DIV11_MODE_TX_1: in     vl_logic;
        FFC_DIV11_MODE_TX_2: in     vl_logic;
        FFC_DIV11_MODE_TX_3: in     vl_logic;
        LDR_CORE2TX_0   : in     vl_logic;
        LDR_CORE2TX_1   : in     vl_logic;
        LDR_CORE2TX_2   : in     vl_logic;
        LDR_CORE2TX_3   : in     vl_logic;
        FFC_LDR_CORE2TX_EN_0: in     vl_logic;
        FFC_LDR_CORE2TX_EN_1: in     vl_logic;
        FFC_LDR_CORE2TX_EN_2: in     vl_logic;
        FFC_LDR_CORE2TX_EN_3: in     vl_logic;
        PCIE_POWERDOWN_0_0: in     vl_logic;
        PCIE_POWERDOWN_0_1: in     vl_logic;
        PCIE_POWERDOWN_1_0: in     vl_logic;
        PCIE_POWERDOWN_1_1: in     vl_logic;
        PCIE_POWERDOWN_2_0: in     vl_logic;
        PCIE_POWERDOWN_2_1: in     vl_logic;
        PCIE_POWERDOWN_3_0: in     vl_logic;
        PCIE_POWERDOWN_3_1: in     vl_logic;
        PCIE_RXPOLARITY_0: in     vl_logic;
        PCIE_RXPOLARITY_1: in     vl_logic;
        PCIE_RXPOLARITY_2: in     vl_logic;
        PCIE_RXPOLARITY_3: in     vl_logic;
        PCIE_TXCOMPLIANCE_0: in     vl_logic;
        PCIE_TXCOMPLIANCE_1: in     vl_logic;
        PCIE_TXCOMPLIANCE_2: in     vl_logic;
        PCIE_TXCOMPLIANCE_3: in     vl_logic;
        PCIE_TXDETRX_PR2TLB_0: in     vl_logic;
        PCIE_TXDETRX_PR2TLB_1: in     vl_logic;
        PCIE_TXDETRX_PR2TLB_2: in     vl_logic;
        PCIE_TXDETRX_PR2TLB_3: in     vl_logic;
        SCIADDR0        : in     vl_logic;
        SCIADDR1        : in     vl_logic;
        SCIADDR2        : in     vl_logic;
        SCIADDR3        : in     vl_logic;
        SCIADDR4        : in     vl_logic;
        SCIADDR5        : in     vl_logic;
        SCIENAUX        : in     vl_logic;
        SCIENCH0        : in     vl_logic;
        SCIENCH1        : in     vl_logic;
        SCIENCH2        : in     vl_logic;
        SCIENCH3        : in     vl_logic;
        SCIRD           : in     vl_logic;
        SCISELAUX       : in     vl_logic;
        SCISELCH0       : in     vl_logic;
        SCISELCH1       : in     vl_logic;
        SCISELCH2       : in     vl_logic;
        SCISELCH3       : in     vl_logic;
        SCIWDATA0       : in     vl_logic;
        SCIWDATA1       : in     vl_logic;
        SCIWDATA2       : in     vl_logic;
        SCIWDATA3       : in     vl_logic;
        SCIWDATA4       : in     vl_logic;
        SCIWDATA5       : in     vl_logic;
        SCIWDATA6       : in     vl_logic;
        SCIWDATA7       : in     vl_logic;
        SCIWSTN         : in     vl_logic;
        HDOUTN0         : out    vl_logic;
        HDOUTN1         : out    vl_logic;
        HDOUTN2         : out    vl_logic;
        HDOUTN3         : out    vl_logic;
        HDOUTP0         : out    vl_logic;
        HDOUTP1         : out    vl_logic;
        HDOUTP2         : out    vl_logic;
        HDOUTP3         : out    vl_logic;
        COUT0           : out    vl_logic;
        COUT1           : out    vl_logic;
        COUT2           : out    vl_logic;
        COUT3           : out    vl_logic;
        COUT4           : out    vl_logic;
        COUT5           : out    vl_logic;
        COUT6           : out    vl_logic;
        COUT7           : out    vl_logic;
        COUT8           : out    vl_logic;
        COUT9           : out    vl_logic;
        COUT10          : out    vl_logic;
        COUT11          : out    vl_logic;
        COUT12          : out    vl_logic;
        COUT13          : out    vl_logic;
        COUT14          : out    vl_logic;
        COUT15          : out    vl_logic;
        COUT16          : out    vl_logic;
        COUT17          : out    vl_logic;
        COUT18          : out    vl_logic;
        COUT19          : out    vl_logic;
        FF_RX_D_0_0     : out    vl_logic;
        FF_RX_D_0_1     : out    vl_logic;
        FF_RX_D_0_2     : out    vl_logic;
        FF_RX_D_0_3     : out    vl_logic;
        FF_RX_D_0_4     : out    vl_logic;
        FF_RX_D_0_5     : out    vl_logic;
        FF_RX_D_0_6     : out    vl_logic;
        FF_RX_D_0_7     : out    vl_logic;
        FF_RX_D_0_8     : out    vl_logic;
        FF_RX_D_0_9     : out    vl_logic;
        FF_RX_D_0_10    : out    vl_logic;
        FF_RX_D_0_11    : out    vl_logic;
        FF_RX_D_0_12    : out    vl_logic;
        FF_RX_D_0_13    : out    vl_logic;
        FF_RX_D_0_14    : out    vl_logic;
        FF_RX_D_0_15    : out    vl_logic;
        FF_RX_D_0_16    : out    vl_logic;
        FF_RX_D_0_17    : out    vl_logic;
        FF_RX_D_0_18    : out    vl_logic;
        FF_RX_D_0_19    : out    vl_logic;
        FF_RX_D_0_20    : out    vl_logic;
        FF_RX_D_0_21    : out    vl_logic;
        FF_RX_D_0_22    : out    vl_logic;
        FF_RX_D_0_23    : out    vl_logic;
        FF_RX_D_1_0     : out    vl_logic;
        FF_RX_D_1_1     : out    vl_logic;
        FF_RX_D_1_2     : out    vl_logic;
        FF_RX_D_1_3     : out    vl_logic;
        FF_RX_D_1_4     : out    vl_logic;
        FF_RX_D_1_5     : out    vl_logic;
        FF_RX_D_1_6     : out    vl_logic;
        FF_RX_D_1_7     : out    vl_logic;
        FF_RX_D_1_8     : out    vl_logic;
        FF_RX_D_1_9     : out    vl_logic;
        FF_RX_D_1_10    : out    vl_logic;
        FF_RX_D_1_11    : out    vl_logic;
        FF_RX_D_1_12    : out    vl_logic;
        FF_RX_D_1_13    : out    vl_logic;
        FF_RX_D_1_14    : out    vl_logic;
        FF_RX_D_1_15    : out    vl_logic;
        FF_RX_D_1_16    : out    vl_logic;
        FF_RX_D_1_17    : out    vl_logic;
        FF_RX_D_1_18    : out    vl_logic;
        FF_RX_D_1_19    : out    vl_logic;
        FF_RX_D_1_20    : out    vl_logic;
        FF_RX_D_1_21    : out    vl_logic;
        FF_RX_D_1_22    : out    vl_logic;
        FF_RX_D_1_23    : out    vl_logic;
        FF_RX_D_2_0     : out    vl_logic;
        FF_RX_D_2_1     : out    vl_logic;
        FF_RX_D_2_2     : out    vl_logic;
        FF_RX_D_2_3     : out    vl_logic;
        FF_RX_D_2_4     : out    vl_logic;
        FF_RX_D_2_5     : out    vl_logic;
        FF_RX_D_2_6     : out    vl_logic;
        FF_RX_D_2_7     : out    vl_logic;
        FF_RX_D_2_8     : out    vl_logic;
        FF_RX_D_2_9     : out    vl_logic;
        FF_RX_D_2_10    : out    vl_logic;
        FF_RX_D_2_11    : out    vl_logic;
        FF_RX_D_2_12    : out    vl_logic;
        FF_RX_D_2_13    : out    vl_logic;
        FF_RX_D_2_14    : out    vl_logic;
        FF_RX_D_2_15    : out    vl_logic;
        FF_RX_D_2_16    : out    vl_logic;
        FF_RX_D_2_17    : out    vl_logic;
        FF_RX_D_2_18    : out    vl_logic;
        FF_RX_D_2_19    : out    vl_logic;
        FF_RX_D_2_20    : out    vl_logic;
        FF_RX_D_2_21    : out    vl_logic;
        FF_RX_D_2_22    : out    vl_logic;
        FF_RX_D_2_23    : out    vl_logic;
        FF_RX_D_3_0     : out    vl_logic;
        FF_RX_D_3_1     : out    vl_logic;
        FF_RX_D_3_2     : out    vl_logic;
        FF_RX_D_3_3     : out    vl_logic;
        FF_RX_D_3_4     : out    vl_logic;
        FF_RX_D_3_5     : out    vl_logic;
        FF_RX_D_3_6     : out    vl_logic;
        FF_RX_D_3_7     : out    vl_logic;
        FF_RX_D_3_8     : out    vl_logic;
        FF_RX_D_3_9     : out    vl_logic;
        FF_RX_D_3_10    : out    vl_logic;
        FF_RX_D_3_11    : out    vl_logic;
        FF_RX_D_3_12    : out    vl_logic;
        FF_RX_D_3_13    : out    vl_logic;
        FF_RX_D_3_14    : out    vl_logic;
        FF_RX_D_3_15    : out    vl_logic;
        FF_RX_D_3_16    : out    vl_logic;
        FF_RX_D_3_17    : out    vl_logic;
        FF_RX_D_3_18    : out    vl_logic;
        FF_RX_D_3_19    : out    vl_logic;
        FF_RX_D_3_20    : out    vl_logic;
        FF_RX_D_3_21    : out    vl_logic;
        FF_RX_D_3_22    : out    vl_logic;
        FF_RX_D_3_23    : out    vl_logic;
        FF_RX_F_CLK_0   : out    vl_logic;
        FF_RX_F_CLK_1   : out    vl_logic;
        FF_RX_F_CLK_2   : out    vl_logic;
        FF_RX_F_CLK_3   : out    vl_logic;
        FF_RX_H_CLK_0   : out    vl_logic;
        FF_RX_H_CLK_1   : out    vl_logic;
        FF_RX_H_CLK_2   : out    vl_logic;
        FF_RX_H_CLK_3   : out    vl_logic;
        FF_TX_F_CLK_0   : out    vl_logic;
        FF_TX_F_CLK_1   : out    vl_logic;
        FF_TX_F_CLK_2   : out    vl_logic;
        FF_TX_F_CLK_3   : out    vl_logic;
        FF_TX_H_CLK_0   : out    vl_logic;
        FF_TX_H_CLK_1   : out    vl_logic;
        FF_TX_H_CLK_2   : out    vl_logic;
        FF_TX_H_CLK_3   : out    vl_logic;
        FFS_CC_OVERRUN_0: out    vl_logic;
        FFS_CC_OVERRUN_1: out    vl_logic;
        FFS_CC_OVERRUN_2: out    vl_logic;
        FFS_CC_OVERRUN_3: out    vl_logic;
        FFS_CC_UNDERRUN_0: out    vl_logic;
        FFS_CC_UNDERRUN_1: out    vl_logic;
        FFS_CC_UNDERRUN_2: out    vl_logic;
        FFS_CC_UNDERRUN_3: out    vl_logic;
        FFS_LS_SYNC_STATUS_0: out    vl_logic;
        FFS_LS_SYNC_STATUS_1: out    vl_logic;
        FFS_LS_SYNC_STATUS_2: out    vl_logic;
        FFS_LS_SYNC_STATUS_3: out    vl_logic;
        FFS_CDR_TRAIN_DONE_0: out    vl_logic;
        FFS_CDR_TRAIN_DONE_1: out    vl_logic;
        FFS_CDR_TRAIN_DONE_2: out    vl_logic;
        FFS_CDR_TRAIN_DONE_3: out    vl_logic;
        FFS_PCIE_CON_0  : out    vl_logic;
        FFS_PCIE_CON_1  : out    vl_logic;
        FFS_PCIE_CON_2  : out    vl_logic;
        FFS_PCIE_CON_3  : out    vl_logic;
        FFS_PCIE_DONE_0 : out    vl_logic;
        FFS_PCIE_DONE_1 : out    vl_logic;
        FFS_PCIE_DONE_2 : out    vl_logic;
        FFS_PCIE_DONE_3 : out    vl_logic;
        FFS_PLOL        : out    vl_logic;
        FFS_RLOL_0      : out    vl_logic;
        FFS_RLOL_1      : out    vl_logic;
        FFS_RLOL_2      : out    vl_logic;
        FFS_RLOL_3      : out    vl_logic;
        FFS_RLOS_HI_0   : out    vl_logic;
        FFS_RLOS_HI_1   : out    vl_logic;
        FFS_RLOS_HI_2   : out    vl_logic;
        FFS_RLOS_HI_3   : out    vl_logic;
        FFS_RLOS_LO_0   : out    vl_logic;
        FFS_RLOS_LO_1   : out    vl_logic;
        FFS_RLOS_LO_2   : out    vl_logic;
        FFS_RLOS_LO_3   : out    vl_logic;
        FFS_RXFBFIFO_ERROR_0: out    vl_logic;
        FFS_RXFBFIFO_ERROR_1: out    vl_logic;
        FFS_RXFBFIFO_ERROR_2: out    vl_logic;
        FFS_RXFBFIFO_ERROR_3: out    vl_logic;
        FFS_TXFBFIFO_ERROR_0: out    vl_logic;
        FFS_TXFBFIFO_ERROR_1: out    vl_logic;
        FFS_TXFBFIFO_ERROR_2: out    vl_logic;
        FFS_TXFBFIFO_ERROR_3: out    vl_logic;
        PCIE_PHYSTATUS_0: out    vl_logic;
        PCIE_PHYSTATUS_1: out    vl_logic;
        PCIE_PHYSTATUS_2: out    vl_logic;
        PCIE_PHYSTATUS_3: out    vl_logic;
        PCIE_RXVALID_0  : out    vl_logic;
        PCIE_RXVALID_1  : out    vl_logic;
        PCIE_RXVALID_2  : out    vl_logic;
        PCIE_RXVALID_3  : out    vl_logic;
        FFS_SKP_ADDED_0 : out    vl_logic;
        FFS_SKP_ADDED_1 : out    vl_logic;
        FFS_SKP_ADDED_2 : out    vl_logic;
        FFS_SKP_ADDED_3 : out    vl_logic;
        FFS_SKP_DELETED_0: out    vl_logic;
        FFS_SKP_DELETED_1: out    vl_logic;
        FFS_SKP_DELETED_2: out    vl_logic;
        FFS_SKP_DELETED_3: out    vl_logic;
        LDR_RX2CORE_0   : out    vl_logic;
        LDR_RX2CORE_1   : out    vl_logic;
        LDR_RX2CORE_2   : out    vl_logic;
        LDR_RX2CORE_3   : out    vl_logic;
        REFCK2CORE      : out    vl_logic;
        SCIINT          : out    vl_logic;
        SCIRDATA0       : out    vl_logic;
        SCIRDATA1       : out    vl_logic;
        SCIRDATA2       : out    vl_logic;
        SCIRDATA3       : out    vl_logic;
        SCIRDATA4       : out    vl_logic;
        SCIRDATA5       : out    vl_logic;
        SCIRDATA6       : out    vl_logic;
        SCIRDATA7       : out    vl_logic;
        REFCLK_FROM_NQ  : in     vl_logic;
        REFCLK_TO_NQ    : out    vl_logic
    );
end PCSD_sim;
