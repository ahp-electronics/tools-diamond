library verilog;
use verilog.vl_types.all;
entity FSCLK_TREE is
    port(
        A               : in     vl_logic;
        Z               : out    vl_logic
    );
end FSCLK_TREE;
