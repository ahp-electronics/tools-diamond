library verilog;
use verilog.vl_types.all;
entity b2_single_ch_serdes is
    generic(
        pd_time         : integer := 10000000;
        lock_step_time  : integer := 1538460;
        ch_id           : integer := 0
    );
    port(
        HDINPi          : in     vl_logic;
        HDINNi          : in     vl_logic;
        rpwdnb          : in     vl_logic;
        tpwdnb          : in     vl_logic;
        mrstb           : in     vl_logic;
        rrst            : in     vl_logic;
        sync            : in     vl_logic;
        tdi             : in     vl_logic_vector(9 downto 0);
        ck3g4tx         : in     vl_logic;
        refck_rx        : in     vl_logic;
        tdrv_dat_sel    : in     vl_logic_vector(1 downto 0);
        bus8bit_sel     : in     vl_logic;
        plb_r2t_en      : in     vl_logic;
        slb_t2r_en      : in     vl_logic;
        slb_r2t_ck_en   : in     vl_logic;
        slb_r2t_d_en    : in     vl_logic;
        slb_eq2t_en     : in     vl_logic;
        bstpadi         : in     vl_logic;
        sentxi          : in     vl_logic;
        senrxi          : in     vl_logic;
        rx_sdi_en       : in     vl_logic;
        rate_mode_rx    : in     vl_logic;
        rate_mode_tx    : in     vl_logic;
        bist_en         : in     vl_logic;
        bist_ch_sel     : in     vl_logic;
        bist_ptn_sel    : in     vl_logic_vector(2 downto 0);
        bist_head_sel   : in     vl_logic_vector(1 downto 0);
        bist_time_sel   : in     vl_logic;
        bist_res_sel    : in     vl_logic_vector(1 downto 0);
        bist_speed_up   : in     vl_logic;
        bstsds_a0       : in     vl_logic;
        lock2ref        : in     vl_logic;
        lock_diff       : in     vl_logic_vector(1 downto 0);
        pci_en          : in     vl_logic;
        pci_ei_en       : in     vl_logic;
        pci_det_ct      : in     vl_logic;
        rate_sel        : in     vl_logic_vector(1 downto 0);
        prem            : in     vl_logic;
        tdrv_pre_set    : in     vl_logic_vector(2 downto 0);
        rxterm_tx       : in     vl_logic_vector(1 downto 0);
        trdv_amp        : in     vl_logic_vector(1 downto 0);
        rterm_rx        : in     vl_logic_vector(1 downto 0);
        losadj          : in     vl_logic_vector(2 downto 0);
        rcv_dcc_en      : in     vl_logic;
        req_en          : in     vl_logic;
        req_lvl_set     : in     vl_logic;
        ser_iset        : in     vl_logic_vector(1 downto 0);
        req_cfg_set     : in     vl_logic_vector(7 downto 0);
        rterm_rxadj     : in     vl_logic_vector(1 downto 0);
        req_i_set       : in     vl_logic_vector(2 downto 0);
        req_pole_adj_en : in     vl_logic;
        pd_i_set        : in     vl_logic_vector(3 downto 0);
        intbiasiset     : in     vl_logic_vector(2 downto 0);
        extbiasiset     : in     vl_logic_vector(2 downto 0);
        cdr_vco_iset    : in     vl_logic_vector(3 downto 0);
        cdr_ctl_a       : in     vl_logic_vector(7 downto 0);
        cdr_ctl_b       : in     vl_logic_vector(7 downto 0);
        cdr_ctl_c       : in     vl_logic_vector(7 downto 0);
        cdr_ctl_d       : in     vl_logic_vector(7 downto 0);
        cdr_ctl_e       : in     vl_logic_vector(7 downto 0);
        cdr_ctl_f       : in     vl_logic_vector(7 downto 0);
        cdr_ctl_g       : in     vl_logic_vector(7 downto 0);
        half_rate_mode  : in     vl_logic;
        HDOUTPi         : out    vl_logic;
        HDOUTNi         : out    vl_logic;
        tcki            : out    vl_logic;
        rcki            : out    vl_logic;
        rdi             : out    vl_logic_vector(9 downto 0);
        pci_det_done    : out    vl_logic;
        pci_connect     : out    vl_logic;
        bsfpadi         : out    vl_logic;
        rloli           : out    vl_logic;
        rlos_lo         : out    vl_logic;
        rlos_hi         : out    vl_logic;
        bist_rpt        : out    vl_logic_vector(7 downto 0)
    );
end b2_single_ch_serdes;
