library verilog;
use verilog.vl_types.all;
entity algn_cascade is
    generic(
        QUAD            : integer := 8;
        GRP             : integer := 4;
        GRP_SEL         : integer := 2;
        CLK_SEL         : integer := 3
    );
    port(
        pcs_rst_n       : in     vl_logic;
        ext_clk_p1_in   : in     vl_logic;
        ext_clk_p2_in   : in     vl_logic;
        ext_done_in     : in     vl_logic;
        quad_clk        : in     vl_logic_vector;
        quad_rst_n      : in     vl_logic_vector;
        quad_start      : in     vl_logic_vector;
        quad_done       : in     vl_logic_vector;
        quad_and_fp1    : in     vl_logic_vector;
        quad_and_fp0    : in     vl_logic_vector;
        quad_or_fp1     : in     vl_logic_vector;
        quad_or_fp0     : in     vl_logic_vector;
        cascade_en_0    : in     vl_logic;
        cascade_en_1    : in     vl_logic;
        cascade_en_2    : in     vl_logic;
        cascade_en_3    : in     vl_logic;
        cascade_en_4    : in     vl_logic;
        cascade_en_5    : in     vl_logic;
        cascade_en_6    : in     vl_logic;
        cascade_en_7    : in     vl_logic;
        grp_sel_0       : in     vl_logic_vector;
        grp_sel_1       : in     vl_logic_vector;
        grp_sel_2       : in     vl_logic_vector;
        grp_sel_3       : in     vl_logic_vector;
        grp_sel_4       : in     vl_logic_vector;
        grp_sel_5       : in     vl_logic_vector;
        grp_sel_6       : in     vl_logic_vector;
        grp_sel_7       : in     vl_logic_vector;
        clk_sel_0       : in     vl_logic_vector;
        clk_sel_1       : in     vl_logic_vector;
        clk_sel_2       : in     vl_logic_vector;
        clk_sel_3       : in     vl_logic_vector;
        ext_algn_en     : in     vl_logic_vector(1 downto 0);
        cascade_ctrl_72 : in     vl_logic_vector(7 downto 2);
        ext_clk_p1_out  : out    vl_logic;
        ext_clk_p2_out  : out    vl_logic;
        ext_done_out    : out    vl_logic;
        grp_clk_p1      : out    vl_logic_vector;
        grp_clk_p2      : out    vl_logic_vector;
        grp_start       : out    vl_logic_vector;
        grp_done        : out    vl_logic_vector;
        grp_deskew_error: out    vl_logic_vector;
        is_slave0_in    : in     vl_logic;
        is_slave1_in    : in     vl_logic;
        is_slave2_in    : in     vl_logic;
        is_slave3_in    : in     vl_logic;
        grp0_wrst_in_n  : in     vl_logic;
        grp1_wrst_in_n  : in     vl_logic;
        grp2_wrst_in_n  : in     vl_logic;
        grp3_wrst_in_n  : in     vl_logic;
        grp0_rrst_in_n  : in     vl_logic;
        grp1_rrst_in_n  : in     vl_logic;
        grp2_rrst_in_n  : in     vl_logic;
        grp3_rrst_in_n  : in     vl_logic;
        is_slave0_out   : out    vl_logic;
        is_slave1_out   : out    vl_logic;
        is_slave2_out   : out    vl_logic;
        is_slave3_out   : out    vl_logic;
        grp0_wrst_out_n : out    vl_logic;
        grp1_wrst_out_n : out    vl_logic;
        grp2_wrst_out_n : out    vl_logic;
        grp3_wrst_out_n : out    vl_logic;
        grp0_rrst_out_n : out    vl_logic;
        grp1_rrst_out_n : out    vl_logic;
        grp2_rrst_out_n : out    vl_logic;
        grp3_rrst_out_n : out    vl_logic
    );
end algn_cascade;
