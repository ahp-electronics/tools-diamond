library verilog;
use verilog.vl_types.all;
entity pcs_channel_top is
    port(
        bus8bit_sel     : in     vl_logic;
        bist_rx_data_sel: in     vl_logic;
        char_mode       : in     vl_logic;
        char_test_data  : in     vl_logic_vector(9 downto 0);
        char_test_mode  : in     vl_logic;
        ebrd_clk        : in     vl_logic;
        fb_clk          : in     vl_logic;
        ff_ebrd_clk     : in     vl_logic;
        ff_rxi_clk      : in     vl_logic;
        ff_tx_d         : in     vl_logic_vector(23 downto 0);
        ff_txi_clk      : in     vl_logic;
        ffc_ei_en       : in     vl_logic;
        ffc_enable_cgalign: in     vl_logic;
        ffc_fb_loopback : in     vl_logic;
        ffc_lane_rx_rst : in     vl_logic;
        ffc_lane_tx_rst : in     vl_logic;
        ffc_pci_det_en  : in     vl_logic;
        ffc_pcie_ct     : in     vl_logic;
        ffc_pfifo_clr   : in     vl_logic;
        ffc_rxpwdnb     : in     vl_logic;
        ffc_rx_div11_clk: in     vl_logic;
        ffc_tx_div11_clk: in     vl_logic;
        ffc_rx_rate_mode: in     vl_logic;
        ffc_tx_rate_mode: in     vl_logic;
        ffc_sb_inv_rx   : in     vl_logic;
        ffc_sb_pfifo_lp : in     vl_logic;
        ffc_signal_detect: in     vl_logic;
        ffc_txpwdnb     : in     vl_logic;
        ffr_clk         : in     vl_logic;
        fft_clk         : in     vl_logic;
        fmbist_data     : in     vl_logic_vector(9 downto 0);
        force_int       : in     vl_logic;
        ion_delay       : in     vl_logic;
        ffc_ldr_core2tx_en: in     vl_logic;
        mc1_chif_ctl    : in     vl_logic_vector(207 downto 0);
        pcie_connect    : in     vl_logic;
        pcie_det_done   : in     vl_logic;
        pcie_powerdown  : in     vl_logic_vector(1 downto 0);
        pcie_rxpolarity : in     vl_logic;
        pcie_txcompliance: in     vl_logic;
        pcie_txdetrx_pr2tlb: in     vl_logic;
        pcie_txelecidle : in     vl_logic;
        pcs_addri       : in     vl_logic_vector(5 downto 0);
        pcs_ctl_3_qd_02 : in     vl_logic_vector(7 downto 0);
        pcs_ctl_4_qd_03 : in     vl_logic_vector(7 downto 0);
        pcs_inti        : in     vl_logic;
        pcs_rdatai      : in     vl_logic_vector(7 downto 0);
        pcs_rdi         : in     vl_logic;
        pcs_wdatai      : in     vl_logic_vector(7 downto 0);
        pcs_wstbi       : in     vl_logic;
        plol            : in     vl_logic;
        quad_reset_all  : in     vl_logic;
        quad_reset_all_n: in     vl_logic;
        rlol            : in     vl_logic;
        rlos_hi         : in     vl_logic;
        rlos_lo         : in     vl_logic;
        rst_ebrd_clk_n  : in     vl_logic;
        rst_fb_clk_n    : in     vl_logic;
        rst_rx_clk_n    : in     vl_logic;
        rst_tx_clk_n    : in     vl_logic;
        rx_clk          : in     vl_logic;
        sci_resetn      : in     vl_logic;
        sciench         : in     vl_logic;
        sciselch        : in     vl_logic;
        sd_rx_clk       : in     vl_logic;
        sd_tx_clk       : in     vl_logic;
        ser_sts_2_ch_27 : in     vl_logic_vector(7 downto 0);
        ser_sts_3_ch_28 : in     vl_logic_vector(7 downto 0);
        ser_sts_4_ch_29 : in     vl_logic_vector(7 downto 0);
        ser_sts_6_ch_2b : in     vl_logic_vector(7 downto 0);
        ser_sts_7_ch_2c : in     vl_logic_vector(7 downto 0);
        serdes_rxd      : in     vl_logic_vector(9 downto 0);
        test_clk        : in     vl_logic;
        tx_clk          : in     vl_logic;
        xge_mode        : in     vl_logic;
        ctie_low        : out    vl_logic;
        ebrd_clk_o      : out    vl_logic;
        fb_clk_o        : out    vl_logic;
        ff_rx_d         : out    vl_logic_vector(23 downto 0);
        ff_rx_f_clk     : out    vl_logic;
        ff_rx_h_clk     : out    vl_logic;
        ff_tx_f_clk     : out    vl_logic;
        ff_tx_h_clk     : out    vl_logic;
        fff_pci_det_en  : out    vl_logic;
        ffr_clk_o       : out    vl_logic;
        ffs_cc_overrun  : out    vl_logic;
        ffs_cc_underrun : out    vl_logic;
        ffs_ls_sync_status: out    vl_logic;
        ffs_rxfbfifo_error: out    vl_logic;
        ffs_txfbfifo_error: out    vl_logic;
        fft_clk_o       : out    vl_logic;
        int_cha_out     : out    vl_logic;
        pcie_beacon_en  : out    vl_logic;
        pcie_mode       : out    vl_logic;
        pcie_phystatus  : out    vl_logic;
        pcie_rxvalid    : out    vl_logic;
        skp_added       : out    vl_logic;
        skp_deleted     : out    vl_logic;
        pcs_addro       : out    vl_logic_vector(5 downto 0);
        pcs_into        : out    vl_logic;
        pcs_rdatao      : out    vl_logic_vector(7 downto 0);
        pcs_rdo         : out    vl_logic;
        pcs_wdatao      : out    vl_logic_vector(7 downto 0);
        pcs_wstbo       : out    vl_logic;
        rst_ebrd_clk_n_o: out    vl_logic;
        rst_fb_clk_n_o  : out    vl_logic;
        rst_rx_clk_n_o  : out    vl_logic;
        rst_tx_clk_n_o  : out    vl_logic;
        rx_ch           : out    vl_logic;
        rx_clk_o        : out    vl_logic;
        sb_txd          : out    vl_logic_vector(9 downto 0);
        ser_ctl_1_ch_10 : out    vl_logic_vector(7 downto 0);
        ser_ctl_2_ch_11 : out    vl_logic_vector(7 downto 0);
        ser_ctl_3_ch_12 : out    vl_logic_vector(7 downto 0);
        ser_ctl_4_ch_13 : out    vl_logic_vector(7 downto 0);
        ser_ctl_5_ch_14 : out    vl_logic_vector(7 downto 0);
        ser_ctl_6_ch_15 : out    vl_logic_vector(7 downto 0);
        ser_ctl_7_ch_16 : out    vl_logic_vector(7 downto 0);
        ser_ch_rst      : out    vl_logic_vector(2 downto 0);
        tobist_data     : out    vl_logic_vector(9 downto 0);
        tsd_pcie_det_ct : out    vl_logic;
        tsd_pcie_ei_en  : out    vl_logic;
        tx_clk_o        : out    vl_logic
    );
end pcs_channel_top;
