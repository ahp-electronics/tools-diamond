library verilog;
use verilog.vl_types.all;
entity I2CA is
    generic(
        I2C_ID          : string  := "I2C0";
        I2C_ADDRESSING  : string  := "7BIT";
        I2C_SLAVE_ADDR  : string  := "0b1000001";
        I2C_BUS_PERF    : string  := "100kHz";
        I2C_CLK_DIVIDER : integer := 1;
        I2C_GEN_CALL    : string  := "DISABLED";
        I2C_INTR_ARBIT  : string  := "DISABLED";
        I2C_INTR_TXRXRDY: string  := "DISABLED";
        I2C_INTR_NACK   : string  := "DISABLED";
        I2C_INTR_GC     : string  := "DISABLED";
        I2C_WAKEUP_SLAVE: string  := "DISABLED";
        I2C_WAKEUP_MASTER: string  := "DISABLED";
        SDA_I_DELAY     : integer := 0;
        SDA_O_DELAY     : integer := 0;
        I2C_FIFO_ENB    : string  := "DISABLED";
        I2C_FIFO_CLKSTR : string  := "DISABLED";
        I2C_FIFO_RXALMOSTF: integer := 30;
        I2C_FIFO_TXALMOSTE: integer := 3;
        I2C_FIFO_INTR_GC: string  := "DISABLED";
        I2C_FIFO_INTR_NACK: string  := "DISABLED";
        I2C_FIFO_MRXRDY : string  := "DISABLED";
        I2C_FIFO_INTR_ARBIT: string  := "DISABLED";
        I2C_FIFO_TXSYNC : string  := "DISABLED";
        I2C_FIFO_TXUNDER: string  := "DISABLED";
        I2C_FIFO_RXOVER : string  := "DISABLED"
    );
    port(
        CSI             : in     vl_logic;
        CLKI            : in     vl_logic;
        STBI            : in     vl_logic;
        WEI             : in     vl_logic;
        ADRI3           : in     vl_logic;
        ADRI2           : in     vl_logic;
        ADRI1           : in     vl_logic;
        ADRI0           : in     vl_logic;
        DATI9           : in     vl_logic;
        DATI8           : in     vl_logic;
        DATI7           : in     vl_logic;
        DATI6           : in     vl_logic;
        DATI5           : in     vl_logic;
        DATI4           : in     vl_logic;
        DATI3           : in     vl_logic;
        DATI2           : in     vl_logic;
        DATI1           : in     vl_logic;
        DATI0           : in     vl_logic;
        DATO9           : out    vl_logic;
        DATO8           : out    vl_logic;
        DATO7           : out    vl_logic;
        DATO6           : out    vl_logic;
        DATO5           : out    vl_logic;
        DATO4           : out    vl_logic;
        DATO3           : out    vl_logic;
        DATO2           : out    vl_logic;
        DATO1           : out    vl_logic;
        DATO0           : out    vl_logic;
        ACKO            : out    vl_logic;
        I2CIRQ          : out    vl_logic;
        I2CWKUP         : out    vl_logic;
        PMUWKUP         : out    vl_logic;
        FIFORST         : in     vl_logic;
        MRDCMPL         : out    vl_logic;
        SRDWR           : out    vl_logic;
        TXFIFOAE        : out    vl_logic;
        TXFIFOE         : out    vl_logic;
        TXFIFOF         : out    vl_logic;
        RXFIFOE         : out    vl_logic;
        RXFIFOAF        : out    vl_logic;
        RXFIFOF         : out    vl_logic;
        SCLI            : in     vl_logic;
        SCLO            : out    vl_logic;
        SCLOEN          : out    vl_logic;
        SDAI            : in     vl_logic;
        SDAO            : out    vl_logic;
        SDAOEN          : out    vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of I2C_ID : constant is 1;
    attribute mti_svvh_generic_type of I2C_ADDRESSING : constant is 1;
    attribute mti_svvh_generic_type of I2C_SLAVE_ADDR : constant is 1;
    attribute mti_svvh_generic_type of I2C_BUS_PERF : constant is 1;
    attribute mti_svvh_generic_type of I2C_CLK_DIVIDER : constant is 1;
    attribute mti_svvh_generic_type of I2C_GEN_CALL : constant is 1;
    attribute mti_svvh_generic_type of I2C_INTR_ARBIT : constant is 1;
    attribute mti_svvh_generic_type of I2C_INTR_TXRXRDY : constant is 1;
    attribute mti_svvh_generic_type of I2C_INTR_NACK : constant is 1;
    attribute mti_svvh_generic_type of I2C_INTR_GC : constant is 1;
    attribute mti_svvh_generic_type of I2C_WAKEUP_SLAVE : constant is 1;
    attribute mti_svvh_generic_type of I2C_WAKEUP_MASTER : constant is 1;
    attribute mti_svvh_generic_type of SDA_I_DELAY : constant is 1;
    attribute mti_svvh_generic_type of SDA_O_DELAY : constant is 1;
    attribute mti_svvh_generic_type of I2C_FIFO_ENB : constant is 1;
    attribute mti_svvh_generic_type of I2C_FIFO_CLKSTR : constant is 1;
    attribute mti_svvh_generic_type of I2C_FIFO_RXALMOSTF : constant is 1;
    attribute mti_svvh_generic_type of I2C_FIFO_TXALMOSTE : constant is 1;
    attribute mti_svvh_generic_type of I2C_FIFO_INTR_GC : constant is 1;
    attribute mti_svvh_generic_type of I2C_FIFO_INTR_NACK : constant is 1;
    attribute mti_svvh_generic_type of I2C_FIFO_MRXRDY : constant is 1;
    attribute mti_svvh_generic_type of I2C_FIFO_INTR_ARBIT : constant is 1;
    attribute mti_svvh_generic_type of I2C_FIFO_TXSYNC : constant is 1;
    attribute mti_svvh_generic_type of I2C_FIFO_TXUNDER : constant is 1;
    attribute mti_svvh_generic_type of I2C_FIFO_RXOVER : constant is 1;
end I2CA;
