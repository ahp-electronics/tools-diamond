library verilog;
use verilog.vl_types.all;
entity b2top_quad is
    port(
        HDINP0          : in     vl_logic;
        HDINN0          : in     vl_logic;
        HDINP1          : in     vl_logic;
        HDINN1          : in     vl_logic;
        HDINP2          : in     vl_logic;
        HDINN2          : in     vl_logic;
        HDINP3          : in     vl_logic;
        HDINN3          : in     vl_logic;
        REFCLKP         : in     vl_logic;
        REFCLKN         : in     vl_logic;
        RXREFCLKP       : in     vl_logic;
        RXREFCLKN       : in     vl_logic;
        ck_core_tx      : in     vl_logic;
        ck_core_rx      : in     vl_logic;
        pwr_on_rst      : in     vl_logic;
        macropdb        : in     vl_logic;
        macrorst        : in     vl_logic;
        trst            : in     vl_logic;
        rrst0           : in     vl_logic;
        rrst1           : in     vl_logic;
        rrst2           : in     vl_logic;
        rrst3           : in     vl_logic;
        td0             : in     vl_logic_vector(9 downto 0);
        td1             : in     vl_logic_vector(9 downto 0);
        td2             : in     vl_logic_vector(9 downto 0);
        td3             : in     vl_logic_vector(9 downto 0);
        rx_sdi_en0      : in     vl_logic;
        rx_sdi_en1      : in     vl_logic;
        rx_sdi_en2      : in     vl_logic;
        rx_sdi_en3      : in     vl_logic;
        pci_en          : in     vl_logic;
        pci_ei_en0      : in     vl_logic;
        pci_ei_en1      : in     vl_logic;
        pci_ei_en2      : in     vl_logic;
        pci_ei_en3      : in     vl_logic;
        pci_det_ct0     : in     vl_logic;
        pci_det_ct1     : in     vl_logic;
        pci_det_ct2     : in     vl_logic;
        pci_det_ct3     : in     vl_logic;
        rpwdnb0         : in     vl_logic;
        rpwdnb1         : in     vl_logic;
        rpwdnb2         : in     vl_logic;
        rpwdnb3         : in     vl_logic;
        tpwdnb0         : in     vl_logic;
        tpwdnb1         : in     vl_logic;
        tpwdnb2         : in     vl_logic;
        tpwdnb3         : in     vl_logic;
        bs2pad_0        : in     vl_logic;
        bs2pad_1        : in     vl_logic;
        bs2pad_2        : in     vl_logic;
        bs2pad_3        : in     vl_logic;
        bstxsel_0       : in     vl_logic;
        bstxsel_1       : in     vl_logic;
        bstxsel_2       : in     vl_logic;
        bstxsel_3       : in     vl_logic;
        bsrxsel_0       : in     vl_logic;
        bsrxsel_1       : in     vl_logic;
        bsrxsel_2       : in     vl_logic;
        bsrxsel_3       : in     vl_logic;
        bsrefclksel     : in     vl_logic;
        bsrxrefclksel   : in     vl_logic;
        rate_sel0       : in     vl_logic_vector(1 downto 0);
        rate_sel1       : in     vl_logic_vector(1 downto 0);
        rate_sel2       : in     vl_logic_vector(1 downto 0);
        rate_sel3       : in     vl_logic_vector(1 downto 0);
        rate_mode_rx0   : in     vl_logic;
        rate_mode_rx1   : in     vl_logic;
        rate_mode_rx2   : in     vl_logic;
        rate_mode_rx3   : in     vl_logic;
        rate_mode_tx0   : in     vl_logic;
        rate_mode_tx1   : in     vl_logic;
        rate_mode_tx2   : in     vl_logic;
        rate_mode_tx3   : in     vl_logic;
        bus8bit_sel     : in     vl_logic;
        tdrv_pre_en0    : in     vl_logic;
        tdrv_pre_en1    : in     vl_logic;
        tdrv_pre_en2    : in     vl_logic;
        tdrv_pre_en3    : in     vl_logic;
        tdrv_pre_set0   : in     vl_logic_vector(2 downto 0);
        tdrv_pre_set1   : in     vl_logic_vector(2 downto 0);
        tdrv_pre_set2   : in     vl_logic_vector(2 downto 0);
        tdrv_pre_set3   : in     vl_logic_vector(2 downto 0);
        rterm_tx0       : in     vl_logic_vector(1 downto 0);
        rterm_tx1       : in     vl_logic_vector(1 downto 0);
        rterm_tx2       : in     vl_logic_vector(1 downto 0);
        rterm_tx3       : in     vl_logic_vector(1 downto 0);
        tdrv_amp0       : in     vl_logic_vector(1 downto 0);
        tdrv_amp1       : in     vl_logic_vector(1 downto 0);
        tdrv_amp2       : in     vl_logic_vector(1 downto 0);
        tdrv_amp3       : in     vl_logic_vector(1 downto 0);
        rterm_rx0       : in     vl_logic_vector(1 downto 0);
        rterm_rx1       : in     vl_logic_vector(1 downto 0);
        rterm_rx2       : in     vl_logic_vector(1 downto 0);
        rterm_rx3       : in     vl_logic_vector(1 downto 0);
        rlos_set        : in     vl_logic_vector(2 downto 0);
        rcv_dcc_en0     : in     vl_logic;
        rcv_dcc_en1     : in     vl_logic;
        rcv_dcc_en2     : in     vl_logic;
        rcv_dcc_en3     : in     vl_logic;
        req_en0         : in     vl_logic;
        req_en1         : in     vl_logic;
        req_en2         : in     vl_logic;
        req_en3         : in     vl_logic;
        req_lvl_set0    : in     vl_logic;
        req_lvl_set1    : in     vl_logic;
        req_lvl_set2    : in     vl_logic;
        req_lvl_set3    : in     vl_logic;
        refck_dcc_en    : in     vl_logic;
        rxrefck_dcc_en  : in     vl_logic;
        refck_core_en   : in     vl_logic;
        rxrefck_en      : in     vl_logic;
        refck_mode      : in     vl_logic_vector(1 downto 0);
        refck_loc_set   : in     vl_logic_vector(1 downto 0);
        refck_rterm     : in     vl_logic;
        tx_ctl_a        : in     vl_logic_vector(7 downto 0);
        tx_ctl_b        : in     vl_logic_vector(7 downto 0);
        tx_ctl_c        : in     vl_logic_vector(7 downto 0);
        tx_ctl_d        : in     vl_logic_vector(7 downto 0);
        rx_ctl_a        : in     vl_logic_vector(7 downto 0);
        rx_ctl_b        : in     vl_logic_vector(7 downto 0);
        rx_ctl_c        : in     vl_logic_vector(7 downto 0);
        rx_ctl_d        : in     vl_logic_vector(7 downto 0);
        rx_ctl_e        : in     vl_logic_vector(7 downto 0);
        rx_ctl_f        : in     vl_logic_vector(7 downto 0);
        rx_ctl_g        : in     vl_logic_vector(7 downto 0);
        rx_ctl_h        : in     vl_logic_vector(7 downto 0);
        cdr_ctl_a0      : in     vl_logic_vector(7 downto 0);
        cdr_ctl_b0      : in     vl_logic_vector(7 downto 0);
        cdr_ctl_c0      : in     vl_logic_vector(7 downto 0);
        cdr_ctl_d0      : in     vl_logic_vector(7 downto 0);
        cdr_ctl_e0      : in     vl_logic_vector(7 downto 0);
        cdr_ctl_f0      : in     vl_logic_vector(7 downto 0);
        cdr_ctl_g0      : in     vl_logic_vector(7 downto 0);
        cdr_ctl_a1      : in     vl_logic_vector(7 downto 0);
        cdr_ctl_b1      : in     vl_logic_vector(7 downto 0);
        cdr_ctl_c1      : in     vl_logic_vector(7 downto 0);
        cdr_ctl_d1      : in     vl_logic_vector(7 downto 0);
        cdr_ctl_e1      : in     vl_logic_vector(7 downto 0);
        cdr_ctl_f1      : in     vl_logic_vector(7 downto 0);
        cdr_ctl_g1      : in     vl_logic_vector(7 downto 0);
        cdr_ctl_a2      : in     vl_logic_vector(7 downto 0);
        cdr_ctl_b2      : in     vl_logic_vector(7 downto 0);
        cdr_ctl_c2      : in     vl_logic_vector(7 downto 0);
        cdr_ctl_d2      : in     vl_logic_vector(7 downto 0);
        cdr_ctl_e2      : in     vl_logic_vector(7 downto 0);
        cdr_ctl_f2      : in     vl_logic_vector(7 downto 0);
        cdr_ctl_g2      : in     vl_logic_vector(7 downto 0);
        cdr_ctl_a3      : in     vl_logic_vector(7 downto 0);
        cdr_ctl_b3      : in     vl_logic_vector(7 downto 0);
        cdr_ctl_c3      : in     vl_logic_vector(7 downto 0);
        cdr_ctl_d3      : in     vl_logic_vector(7 downto 0);
        cdr_ctl_e3      : in     vl_logic_vector(7 downto 0);
        cdr_ctl_f3      : in     vl_logic_vector(7 downto 0);
        cdr_ctl_g3      : in     vl_logic_vector(7 downto 0);
        pll_ctl_a       : in     vl_logic_vector(7 downto 0);
        pll_ctl_b       : in     vl_logic_vector(7 downto 0);
        pll_ctl_c       : in     vl_logic_vector(7 downto 0);
        pll_ctl_d       : in     vl_logic_vector(7 downto 0);
        pll_ctl_e       : in     vl_logic_vector(7 downto 0);
        pll_ctl_f       : in     vl_logic_vector(7 downto 0);
        pll_ctl_g       : in     vl_logic_vector(7 downto 0);
        ibias_a         : in     vl_logic_vector(7 downto 0);
        bstsds_a        : in     vl_logic_vector(7 downto 0);
        bstsds_b        : in     vl_logic_vector(7 downto 0);
        bstsds_c        : in     vl_logic_vector(7 downto 0);
        RESP            : inout  vl_logic;
        VDDIB0          : in     vl_logic;
        VDDIB1          : in     vl_logic;
        VDDIB2          : in     vl_logic;
        VDDIB3          : in     vl_logic;
        VDDOB0          : in     vl_logic;
        VDDOB1          : in     vl_logic;
        VDDOB2          : in     vl_logic;
        VDDOB3          : in     vl_logic;
        VDDAX25         : in     vl_logic;
        VDDRX0          : in     vl_logic;
        VDDRX1          : in     vl_logic;
        VDDRX2          : in     vl_logic;
        VDDRX3          : in     vl_logic;
        VDDTX0          : in     vl_logic;
        VDDTX1          : in     vl_logic;
        VDDTX2          : in     vl_logic;
        VDDTX3          : in     vl_logic;
        VSSRX           : in     vl_logic;
        VSSTX           : in     vl_logic;
        VDDP            : in     vl_logic;
        VSSP            : in     vl_logic;
        iref50_ext_0    : inout  vl_logic;
        iref50_ext_1    : inout  vl_logic;
        iref50_ext_2    : inout  vl_logic;
        iref50_ext_3    : inout  vl_logic;
        iref50_int_0    : inout  vl_logic;
        iref50_int_1    : inout  vl_logic;
        iref50_int_2    : inout  vl_logic;
        iref50_int_3    : inout  vl_logic;
        iref50_ext_in   : inout  vl_logic;
        iref50_int_in   : inout  vl_logic;
        resp_use        : in     vl_logic;
        logic_hi        : out    vl_logic;
        logic_low       : out    vl_logic;
        HDOUTP0         : out    vl_logic;
        HDOUTN0         : out    vl_logic;
        HDOUTP1         : out    vl_logic;
        HDOUTN1         : out    vl_logic;
        HDOUTP2         : out    vl_logic;
        HDOUTN2         : out    vl_logic;
        HDOUTP3         : out    vl_logic;
        HDOUTN3         : out    vl_logic;
        rd0             : out    vl_logic_vector(9 downto 0);
        rd1             : out    vl_logic_vector(9 downto 0);
        rd2             : out    vl_logic_vector(9 downto 0);
        rd3             : out    vl_logic_vector(9 downto 0);
        rck0            : out    vl_logic;
        rck1            : out    vl_logic;
        rck2            : out    vl_logic;
        rck3            : out    vl_logic;
        rlol0           : out    vl_logic;
        rlol1           : out    vl_logic;
        rlol2           : out    vl_logic;
        rlol3           : out    vl_logic;
        rlos_lo0        : out    vl_logic;
        rlos_lo1        : out    vl_logic;
        rlos_lo2        : out    vl_logic;
        rlos_lo3        : out    vl_logic;
        rlos_hi0        : out    vl_logic;
        rlos_hi1        : out    vl_logic;
        rlos_hi2        : out    vl_logic;
        rlos_hi3        : out    vl_logic;
        pci_connect0    : out    vl_logic;
        pci_connect1    : out    vl_logic;
        pci_connect2    : out    vl_logic;
        pci_connect3    : out    vl_logic;
        pci_det_done0   : out    vl_logic;
        pci_det_done1   : out    vl_logic;
        pci_det_done2   : out    vl_logic;
        pci_det_done3   : out    vl_logic;
        tck0            : out    vl_logic;
        tck1            : out    vl_logic;
        tck2            : out    vl_logic;
        tck3            : out    vl_logic;
        refck2core      : out    vl_logic;
        rxrefck2core    : out    vl_logic;
        plol            : out    vl_logic;
        refloc          : out    vl_logic;
        rrefloc         : out    vl_logic;
        bstsds_rpt      : out    vl_logic_vector(7 downto 0);
        bs4pad_0        : out    vl_logic;
        bs4pad_1        : out    vl_logic;
        bs4pad_2        : out    vl_logic;
        bs4pad_3        : out    vl_logic;
        bs4refck        : out    vl_logic;
        bs4rxrefck      : out    vl_logic;
        sds_test_bus    : out    vl_logic_vector(7 downto 0)
    );
end b2top_quad;
