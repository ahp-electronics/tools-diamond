library verilog;
use verilog.vl_types.all;
entity pfalu is
    port(
        clk             : in     vl_logic;
        rst             : in     vl_logic;
        rst_int         : in     vl_logic;
        alu_ok          : in     vl_logic;
        mul_b_adr       : in     vl_logic_vector(8 downto 0);
        alu_a_adr       : in     vl_logic_vector(8 downto 0);
        alu_b_adr       : in     vl_logic_vector(8 downto 0);
        mul_s_adr       : in     vl_logic_vector(8 downto 0);
        mul_s_wr        : in     vl_logic;
        alu_s_adr       : in     vl_logic_vector(8 downto 0);
        alu_s_wr        : in     vl_logic;
        glb_w_adr       : in     vl_logic_vector(8 downto 0);
        glb_w_data      : in     vl_logic_vector(31 downto 0);
        glb_w_wr        : in     vl_logic;
        glb_r_adr2      : in     vl_logic_vector(8 downto 0);
        glb_r_data2     : out    vl_logic_vector(31 downto 0);
        do_sub          : in     vl_logic;
        do_xor          : in     vl_logic;
        do_add          : in     vl_logic;
        do_set          : in     vl_logic;
        do_chk          : in     vl_logic;
        do_mov          : in     vl_logic;
        do_sft1         : in     vl_logic;
        do_sft8         : in     vl_logic;
        do_sft24        : in     vl_logic;
        do_msk          : in     vl_logic;
        do_mul          : in     vl_logic;
        msk_op          : in     vl_logic_vector(1 downto 0);
        msk_set         : in     vl_logic_vector(9 downto 0);
        msk_idx         : in     vl_logic_vector(4 downto 0);
        chk_op          : in     vl_logic;
        use_carry       : in     vl_logic;
        clear_eq        : in     vl_logic;
        sign_ext        : in     vl_logic;
        alu_a_rnd       : in     vl_logic;
        alu_a_36        : in     vl_logic;
        alu_a_5c        : in     vl_logic;
        alu_a_is0       : in     vl_logic;
        alu_a_is1       : in     vl_logic;
        alu_b_sel_u     : in     vl_logic;
        alu_b_ovr       : in     vl_logic;
        alu_co          : out    vl_logic;
        alu_bs          : out    vl_logic;
        alu_sn          : out    vl_logic;
        alu_od          : out    vl_logic;
        alu_eq          : out    vl_logic
    );
end pfalu;
