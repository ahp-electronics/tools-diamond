library verilog;
use verilog.vl_types.all;
entity SLRST_N_TREE is
    port(
        A               : in     vl_logic;
        Z               : out    vl_logic
    );
end SLRST_N_TREE;
