------------------------------------------------------------------------
@E
---a-RERH#VCHDR#ENRR0FL#CREbHbCC8RM$Osb80C!
!!-a-RERH#VCHDRF#EkRD8MCCPsCRLRH#Eb8bCRRHMs8CNNCLDRsVFl!!!

---a-RERH#P#CsHRFMF0VREvCRq_a])p qRObN	CNoR
H#-1-RbHCOVRHO01FR$DMbHRV$NRM8HM#RFk0R#DNLCFRVsHR#lNkD0MHF
R--B$FbsEHo0OR52gR4gRc,1b$MDHHO0R$,Q3MORDqDRosHER0#sCC#s8PC

---a-RE=CR>bRFC0sNFHsR##RkC08RFbR#CVOH$RRNLDkH0MRHRbHlDCClM00NHRFM
R--VRFsN$R0bFCRskRVMHO0F
M3---
-ERaCsRF8RCsFVVRk0MOH#FMR8NMRO8CDNNs0MHF##RHR0MFRCH8MO0HN0DRFER0C-
-RHFsoNHMDCRPsF#HMFRVsCR#OHks0s$RCFN#M
#3---
-]RfCCN8s/:R/M#$bODHH/0$ObFl.jj.j$d#M/b.ObFlHsDC#E/P8PD/El8/N_0EsDCN38PEyf4R

---w-RFwsRkEs0C8sRCs#OHHb0F8MRCH0NDR#,bNDC#DCRFRF	NO0RFCllMR0#LFCDI-:
---------------------------------------------------------------------
-----
-FRBbH$soRE04nggRRL$Q   3DRqDHRso#E0R#sCCCsP8-3
--
-RHaE#FR#kCsORDVHC#RHRRNMCC##MN0HDNRbsF0RV RQ 1 R048Rj3(n.g-4gRn,Q   RN10Ms8N8-R
-]Re7vpRNC0ElHN0ORNDu	NON#oC3ERaH##RFOksCHRVDlCRNM$RFL0RCFROb8HC,FR#DR8,F
sR-H-RMkOD8RC8IEH0RV#F0sINCER0NH0R#FR#DI8RHF0EkI0Rs0H0CbMRCHsl#F#HMsRVF0lREQCR 
  -1-R08NMN#s8Rb7CNls0C3M0RHaE#FR#kCsORDVHCNRl$CRLRCk#8FR0RbHlDCClM00RERH##M0N88NsR-
-R8NMR$lNRRLC80H#skHL0RC8HOMRFHlbDRC8VlFsRRHMNRM$lMNMC#sRFFRDMNoR#ER0C-R
-FROlDbHCV8RFRsl8#FCR0MFRDNDF8IRHOsC0CR8ObFlH0DNHRFMF0VREFCRsHHoMRND#sFkOVCRH3DC
R--a#EHRk#FsROCVCHDR$lNRRLCOHFbCV8RFHsRMP8HHN8kD#RkCCRL0CICMHRDO#CMCk8R##Cs3-R
-ERaH##RFOksCHRVDHCR#sRbF8PHCF8RMMRNRRq1QL1RN##H3ERaC RQ 8 RHD#ON#HlRYqhR-
-R)Wq)aqhYXR u1) 1)RmRuQvp7Q RBQhpQz7hqtRhWYRqq))hRaYmvwR ])BqqhaAQQpa
YR-q-Rhw7RQ ah1w1Rmz)R1w Rmq)RR)uqazQBpRq)uuz)m31 RCaERCk#sVRFRC0ERk#FsROC
R--VCHDRN#EDHDRMl8CM$HVR8NMRDEF8 RQ E RNDslCR##VlsFR$NMRl8NN#oCRRFsDLHNH0DH$-R
-sRNHM#HokRF0VRFRC0ERCk#RC0EsVCF3-
-
R--aDH0CR:RRRRRRN10Ms8N8]Re7vpRNC0ElHN0ORNDu	NON#oCR 5Q 1 R048Rj3(n.g-4gRn,
R--RRRRRRRRRRRRRavq] _)q
p2---
-HRpLssN$R:RRaRRERH#b	NONRoC#DENDCRLRlOFbCHD8MRH0NFRRLDHs$Ns
R--RRRRRRRRRRRRRl#$LHFDODND$NRMlRC8Q   3-
-
R--7CCPDCFbsR#:R Q  qR71eBR]R7pvEN0C0lNHDONROuN	CNo#FRWsM	HosRtF
kb---
-kRus#bFCR:RRaRRERH#b	NONRoC8HCVMRC#N0R#NNM8sV8RF8sRCo#HM#CsRR0FkR#CH-M
-RRRRRRRRRRRR8RRCs#OHMLHo]Re7lpRFD8C#ER0Nl0RNR	CkR#CFOVRFFllM R)qOpRF0M#N#M0
R--RRRRRRRRRRRRR8NMRlOFlRFM)p qRCCDl0CMNRs$lEN0C0lNHDONRMVkOF0HM
#3---
-HRplNH00MHF:aRREPCRNCDk#CRoMNCs0RC8L0$REVCRk0MOH#FMRRHM0#EHRObN	CNoR$lN
R--RRRRRRRRRRRRRsPN$sRVFblRDVN0FRsl0bFRDVN0F,slR8NMRC0ERCbsOHH#FFMRVCRs#0kD#-
-RRRRRRRRRRRRR#RHRDFM$kRoNMsN08CCRR0FL0CRElCRHlMHkslRCHJksRC8LQ$R R  1R084nj(--
-RRRRRRRRRRRRRgR4g
d3---
-FRh0:C#
R--RRRRRRRRRRRRRRhF8DCON0sNH#FMRRFs8HCVMHH0FRM##DENDCRLROHMDCk88MRH,sRF
R--RRRRRRRRRRRRROCGDCk88sRVFRl,0#EHRObN	CNo3-
-RRRRRRRRRRRRRERaCbR"NNO	o8CRCNODsHN0FRM"8HCVMRC#0REC0C$b##,Rk$L0b,C#R8NM
R--RRRRRRRRRRRRRO8CDNNs0MHF#VRFRavq] _)q
p3-R-RRRRRRRRRRRRRaREC#M0N88NsR0lNENCl0NHODCR8VHHM0MHFR8NMRMOFP0CMHNFMDCRlNMMHo-
-RRRRRRRRRRRRRVRFRC0ER0lNENCl0NHODkRVMHO0FRM#00ENRCNsRsbN0VRFRH0E#0R#NNM8s-8
-RRRRRRRRRRRRsRRCCbs#0CMRC0ERsVFlRND#NClMO0H#VRFRC0ERbHlDCClM00NHRFMF0VRE-C
-RRRRRRRRRRRRvRRq_a])p qRObN	CNoRO8CDNNs0MHF3aRREbCRkFsb#FCRVER0CqRva)]_ 
qp-R-RRRRRRRRRRRRRb	NONRoCL$F8RRH#0bFRsHFP8NCRRHok8HCDMVCRFHsRlCbDl0CMNF0HM0#RF-
-RRRRRRRRRRRRRCRPs$HVRC0EHHsRlCbDl0CMNF0HMVRFRavq] _)qRp3RFaFDCR8PFCDb#CsR$lN
R--RRRRRRRRRRRRRFOEFR#C0HFRlCbDl0CMRC0ERObN	CNoR8LF$MRHRC0ER#lF0VRCVHHOC
M0-R-RRRRRRRRRRRRRlMNMCNsRPDNHNCLDRR0F0lEC3-
-
R--------------------------------------------------------------------------------
-RseC#MHFRRRR:3R46-
-R07NCRRRRRRR:cR.RDKk$gR4g-n
--R--------------------------------------------------------------------------
--
#--$EM0C##HR0HMCNsMDN_bOo	NCN
bOo	NCqRva)]_ RqpHR#
RORRF0M#NRM0B$Fb)EHo00hFH:OCR)1aQ
htRRRRR=R:RF"BbH$soRE04nggR Q  q3RDsDRH0oE#CRs#PCsC"83;R

R-RR-R
RR-R-RMBF#M0N0CR7VHHM0MHF#R
RR-R-
RRRRMOF#M0N0vRRq_a]4e_m  )_R):R Rqp:j=R3(dnUg(_c4c4_c(4cd._.j4n;R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-e-RNCDkRRFV4
/CRRRRO#FM00NMRqRva ]_R):R Rqp:.=R3U(4.4U_Uc.U_j6gc.6_dn6d;R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-e-RNCDkRRFVCR
RRFROMN#0MR0Rv]qa_u._QRR:)p qRR:=nU3.d_4U6(dj4g_(6_Uncg(ndR;
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--ekNDCVRFRb.*HR
RRFROMN#0MR0Rv]qa_RuQ: R)q:pR=3Rd46c4gn_.6_d6Ugg(dd_.U;cn
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-NReDRkCFbVRHR
RRFROMN#0MR0Rv]qa__uQm)e _:.RRq) p=R:R643(gj(_.ndng(_cnUg_gn4.
d;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RDeNkFCRVHRb/R.
RORRF0M#NRM0Ravq]__4m)e _RuQ: R)q:pR=3Rjdd4UjU_gU_n4Ugd(j(_n4;6c
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-NReDRkCF4VR/
bHRRRRO#FM00NMRqRvau]_Qe_m d)_R):R Rqp:4=R3(jc4(g_6464_6gng((_c6n4;R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-e-RNCDkRRFVbdH/
RRRRMOF#M0N0vRRq_a]umQ_e_ )cRR:)p qRR:=jU3(6_dgUd4nd(_gc_cUdnjg.R;
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--ekNDCVRFR/bHcR
RRFROMN#0MR0Rv]qa_ud_Qe_m .)_R):R Rqp:c=R3.(4dUU_gdUj_nUcUUg_6g(n;R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-e-RNCDkRbd*H
/.RRRRO#FM00NMRqRvap]_mmt_wR_.: R)q:pR=3Rjn4gdc4_(U_j66cgg6j_dg;c.
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-NRh0NksDFRDoVRFRR.
RORRF0M#NRM0Ravq]m_ptw_m_R4j: R)q:pR=3R.d6j.Uj_6g_.ggccj6U_nc;j.
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-NRh0NksDFRDoVRFR
4jRRRRO#FM00NMRqRvap]_m_t.m w_R):R Rqp:4=R3.ccn6g_jUcj_gUUncd_j;(c
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-FRpoNRL#.CRRRFVCR
RRFROMN#0MR0Rv]qa_tpm4mj_w:_ Rq) p=R:Rcj3dgc._Ucc4jg_d4.6_(U.n
6;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RopFR#LNCjR4RRFVCR
RRFROMN#0MR0Rv]qa_m4_e_ )1aT)_R.:)p qRR:=jj3((_4jn4(U4n_U6_c(6c.cjR;
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--#NJkssCRFRF0F4VR/R.
RORRF0M#NRM0Ravq]T_1).a_: R)q:pR=3R4c.4c46_dn_.d(gdj6c_jU;Uj
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-JR#kCNsRFsF0VRFRR.
RORRF0M#NRM0Ravq] _7tm_a_7)q: R)q:pR=3Rjjc4(6._dg_.64cggdg_.6;((
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RMBFP#CsHRFMV0NOFVsRsRFl8sCoC0CRFNRs8MHN
RRRRMOF#M0N0vRRq_a]1aT)_:uQRq) p=R:R(43(6.c_6dUjjg_6n64_(j.d
j;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-Rk#JNRsCs0FFRRFVbRH
RORRF0M#NRM0Ravq]q_)7m_a_t7 : R)q:pR=(R636.g(g(_6j4d_dU..Uj_(jnU;R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-FRBMsPC#MHFROVN0RFsVlsFR8sNHRNM08FRCCosCR

R-RR-R
RR-R-RMwkOF0HMCR7OsDNNF0HMR#
R-RR-R
RRkRVMHO0FBMR RQp5:XRRRHM)p qRs2RCs0kM R)q
p;RRRRRRRR-u-RkFsb#
C:RRRRRRRR-R-RRRRRR)RRCs0kM##RlDNDCR#0Q hatR )PkNDCNR5# R)qRp2MRF0D#C#RN0EM
RXRRRRRRRR-1-RbHCONPDRNCDk#R:
RRRRR-RR-RRRRRRRRFRhMRC
RRRRR-RR-FR7lMNH:R
RRRRRR-R-RRRRRRRRRHXRM R)qRp
RRRRR-RR-sR sRFsO8FMHF0HM
#:RRRRRRRR-R-RRRRRRhRRF
MCRRRRRRRR-)-RNCMo:R
RRRRRR-R-RRRRRRRRRQB p25XRRH#lEN0C0lNHDONDk$RMkLFM88C
RRRRRRRRR--hCF0#R:
RRRRR-RR-RRRRRRRR2RNRbQlDCClM00NH#FMRPENCFR0Rb#kb0FsRRN0D#CN0ER0CFR8lMNH
RRRRRRRRR--RRRRRRRRRRRRRqRRAX152RR<)p q5aQh )t 't]Q]
2
RRRRVOkM0MHFRt1QhXR5:MRHRq) pRR2skC0s)MR ;qp
RRRRRRRRR--ubksF:#C
RRRRRRRRR--RRRRRRRR)kC0sRM#4R3jHXVRRj>R3Rj;jR3jHXVRRj=R3Rj;-j43RRHVXRR<j
3jRRRRRRRR-1-RbHCONPDRNCDk#R:
RRRRR-RR-RRRRRRRRFRhMRC
RRRRR-RR-FR7lMNH:R
RRRRRR-R-RRRRRRRRRHXRM R)qRp
RRRRR-RR-sR sRFsO8FMHF0HM
#:RRRRRRRR-R-RRRRRRhRRF
MCRRRRRRRR-)-RNCMo:R
RRRRRR-R-RRRRRRRRR1qA5t1Qh25X2=R<Rj43
RRRRRRRRR--hCF0#R:
RRRRR-RR-RRRRRRRRFRhM
C
RRRRVOkM0MHFRz)mh57RXRR:H)MR Rqp2CRs0MksRq) pR;
RRRRR-RR-kRus#bFCR:
RRRRR-RR-RRRRRRRRFR)k#M8R0XRFER0CCRMN#sC0MRH0CCosNRPDRkC5RN#sDCN2Q3RVRRXHR#
RRRRR-RR-RRRRRRRRNREDNVI$CRL0CICMIR0FMRH0CCosR#,sMFk8oHMRRH#N$INRFVsl3RjjR
RRRRRR-R-RC1bODHNRDPNk:C#
RRRRRRRRR--RRRRRRRR)hmz735jj=2RRjj3
RRRRRRRRR--7NFlH
M:RRRRRRRR-R-RRRRRRXRRRRHM)p q
RRRRRRRRR-- FsssFROM08HH#FM:R
RRRRRR-R-RRRRRRRRRMhFCR
RRRRRR-R-RM)No
C:RRRRRRRR-R-RRRRRR)RRm7zh5RX2Hl#RNC0ElHN0ODND$MRkLMFk8
C8RRRRRRRR-h-RF#0C:R
RRRRRR-R-RRRRRRRRRRN2QDlbCMlC0HN0FRM#ECNPRR0F#bkbFRs0ND0RC0N#RC0ERl8FN
HMRRRRRRRR-R-RRRRRRRRRRRRRRARq125XR)<R 5qpQ hat' )]]Qt2R

RVRRk0MOHRFM)p qvRQh5RX,YRR:H)MR Rqp2CRs0MksRq) pR;
RRRRR-RR-kRus#bFCR:
RRRRR-RR-RRRRRRRRCR)0Mks#ER0CDRNosCLNNHODRD$#DlNDRCsFXVRR8NMRRY
RRRRR-RR-bR1CNOHDNRPD#kC:R
RRRRRR-R-RRRRRRRRRq) phvQ5YX,2RR=XERICXMRRY=R
RRRRRRRRR--7NFlH
M:RRRRRRRR-R-RRRRRRXRRRRHM)p q;RRYH)MR 
qpRRRRRRRR- -RsssFRMOF8HH0F:M#
RRRRRRRRR--RRRRRRRRhCFM
RRRRRRRRR--)oNMCR:
RRRRR-RR-RRRRRRRR R)qQpvh,5XYH2R#NRl0lECNO0HN$DDRLkMF8kMCR8
RRRRR-RR-FRh0:C#
RRRRRRRRR--RRRRRRRRhCFM
R
RRkRVMHO0FaMR)BzhRR5X:MRHRq) pRR2skC0s)MR ;qp
RRRRRRRRR--ubksF:#C
RRRRRRRRR--RRRRRRRRaMskOCN0#RRX0NFIsR8#jR3jNRM8skC0sRM#0MskOCN08NRPD
kCRRRRRRRR-1-RbHCONPDRNCDk#R:
RRRRR-RR-RRRRRRRR)Raz5hBj23jRj=R3Rj
RRRRR-RR-FR7lMNH:R
RRRRRR-R-RRRRRRRRRHXRM R)qRp
RRRRR-RR-sR sRFsO8FMHF0HM
#:RRRRRRRR-R-RRRRRRhRRF
MCRRRRRRRR-)-RNCMo:R
RRRRRR-R-RRRRRRRRRza)hXB52#RHR0lNENCl0NHODRD$kFMLkCM88R
RRRRRR-R-R0hFC
#:RRRRRRRR-R-RRRRRRNRR2lRQblDCCNM00MHF#NREP0CRFkR#bsbF00RNRNDC#00RE8CRFHlNMR
RRRRRR-R-RRRRRRRRRRRRRRRRq5A1X<2RRq) ph5Qa  t)Q']t
]2
RRRRMVkOF0HMpRwmRm)5:XRRRHM)p qRs2RCs0kM R)q
p;RRRRRRRR-u-RkFsb#
C:RRRRRRRR-R-RRRRRR)RRCs0kMD#RNCso#Q0Rhta  P)RNCDkR#5NRq) pM2RFo0Rs0CNC0sRERNMXR
RRRRRR-R-RC1bODHNRDPNk:C#
RRRRRRRRR--RRRRRRRRwmpm)35jj=2RRjj3
RRRRRRRRR--7NFlH
M:RRRRRRRR-R-RRRRRRXRRRRHM)p q
RRRRRRRRR-- FsssFROM08HH#FM:R
RRRRRR-R-RRRRRRRRRMhFCR
RRRRRR-R-RM)No
C:RRRRRRRR-R-RRRRRRwRRp)mm5RX2Hl#RNC0ElHN0ODND$MRkLMFk8
C8RRRRRRRR-h-RF#0C:R
RRRRRR-R-RRRRRRRRRRN2QDlbCMlC0HN0FRM#ECNPRR0F#bkbFRs0ND0RC0N#RC0ERl8FN
HMRRRRRRRR-R-RRRRRRRRRRRRRRARq125XR)<R 5qpQ hat' )]]Qt2R

RVRRk0MOHRFM"7vm"XR5,:RYRRHM)p qRs2RCs0kM R)q
p;RRRRRRRR-u-RkFsb#
C:RRRRRRRR-R-RRRRRR)RRCs0kMV#RD0FNHRMobMFH0FRl8kkD#VRFRYX/,HRI00ERE#CRNRlC#MHoR
N#RRRRRRRR-R-RRRRRRYRR,MRN8LRN#kFD0PCRNCDkR#DC#ER0N0MRENCRLD#FkR0CPkNDCVRFRRY,N
M8RRRRRRRR-R-RRRRRRVRRF#sRFRlCQ hatR )PkNDCRRh0RECskC#D#0RN#0HV#HCRC0ERDsCNF0HMR
RRRRRR-R-RRRRRRRRR=XRRhY*Rv+RmX75,
Y2RRRRRRRR-1-RbHCONPDRNCDk#R:
RRRRR-RR-RRRRRRRRFRhMRC
RRRRR-RR-FR7lMNH:R
RRRRRR-R-RRRRRRRRRHXRM R)qRp;YMRHRq) pMRN8RRY/j=R3Rj
RRRRR-RR-sR sRFsO8FMHF0HM
#:RRRRRRRR-R-RRRRRR RRsssFRRHVYRR=j
3jRRRRRRRR-)-RNCMo:R
RRRRRR-R-RRRRRRRRR1qA57vm5YX,2<2RR1qA5
Y2RRRRRRRR-h-RF#0C:R
RRRRRR-R-RRRRRRRRRMhFCR

RVRRk0MOHRFM)p qvRqX5RX,YRR:H)MR Rqp2CRs0MksRq) pR;
RRRRR-RR-kRus#bFCR:
RRRRR-RR-RRRRRRRRCR)0Mks#ER0CDRNosCLNNHODRD$DoNsCFsRVRRXNRM8YR
RRRRRR-R-RC1bODHNRDPNk:C#
RRRRRRRRR--RRRRRRRR)p qv5qXX2,YRX=RRCIEMRRX=
RYRRRRRRRR-7-RFHlNMR:
RRRRR-RR-RRRRRRRRRRXH)MR ;qpRHYRM R)qRp
RRRRR-RR-sR sRFsO8FMHF0HM
#:RRRRRRRR-R-RRRRRRhRRF
MCRRRRRRRR-)-RNCMo:R
RRRRRR-R-RRRRRRRRRq) pXvq5YX,2#RHR0lNENCl0NHODRD$kFMLkCM88R
RRRRRR-R-R0hFC
#:RRRRRRRR-R-RRRRRRhRRF
MC
RRRRMVkOF0HMTR1)5aRXRR:H)MR Rqp2CRs0MksRq) pR;
RRRRR-RR-kRus#bFCR:
RRRRR-RR-RRRRRRRRCR)0Mks#JR#kCNsRFsF0VRFRRX
RRRRR-RR-bR1CNOHDNRPD#kC:R
RRRRRR-R-RRRRRRRRR)1Ta35jj=2RRjj3
RRRRRRRRR--RRRRRRRR1aT)5j432RR=4
3jRRRRRRRR-7-RFHlNMR:
RRRRR-RR-RRRRRRRRRRX>j=R3Rj
RRRRR-RR-sR sRFsO8FMHF0HM
#:RRRRRRRR-R-RRRRRR RRsssFRRHVXRR<j
3jRRRRRRRR-)-RNCMo:R
RRRRRR-R-RRRRRRRRR)1Ta25XRR>=j
3jRRRRRRRR-h-RF#0C:R
RRRRRR-R-RRRRRRRRRRN2aRECkCbbsFRLkRM8F0VREsCRCENONCLDRMsNoFCRVTR1)HaR#R
RRRRRR-R-RRRRRRRRRRRRNsbbFlGHND0C$HRoPRCML
$:RRRRRRRR-R-RRRRRRRRRRRRRRTR1)Xa52=R<R)1Ta 5)q]p'Q2t]
R
RRsRbF8OCkRsCzwhQm5)vPHNsNCLDR 1 714, . 7:FHMku0Rma1QQ;e RsPNHDNLC:RXFRk0)p q2R;
RRRRR-RR-kRus#bFCR:
RRRRR-RR-RRRRRRRRCR)0Mks#H,RM,RXRbNR#8CkFN-sMl8FRlMkLRCsIEH0RHkMVlFs
RRRRRRRRR--RRRRRRRR80H#skHL0MHFRRHM0RECFMbCR0HMCNsPDjR53Rj,423j3R
RRRRRR-R-RC1bODHNRDPNk:C#
RRRRRRRRR--RRRRRRRRhCFM
RRRRRRRRR--7NFlH
M:RRRRRRRR-R-RRRRRR4RRRR<=17  4=R<Rc.4(dcU6;n.R<4R= R1 R7.<.=R4cc(UgddUR
RRRRRR-R-Rs sFOsRFHM80MHF#R:
RRRRR-RR-RRRRRRRRsR sRFsH1VR 4 7RRFs17  .kRF08#HCVRFRDPNH88RFHlNMR
RRRRRR-R-RM)No
C:RRRRRRRR-R-RRRRRRjRR3<jRR<XRRj43
RRRRRRRRR--hCF0#R:
RRRRR-RR-RRRRRRRR2RNRCaERl#CNHM0OV#RF0sRERH#VOkM0MHFRCNsR#8COLsHCL8R$ER0CR
RRRRRR-R-RRRRRRRRRRRRNFDosEH0lkRbL#DHERC8Lu$RHsCsC'Rp $OkCHsRMBR"FkllMNHO0MHF#R
RRRRRR-R-RRRRRRRRRRRRF0VREqCRB"v,RDPF34Rd,FRM3,RnRMKkCgR4URU,bRb3(-c.(3(c
RRRRRRRRR--RRRRRRRRRaRRENCRDsoFHl0ERRH#LCN#8MRFRC0ERlOFLNHM0MHFRRFV0
IFRRRRRRRR-R-RRRRRRRRRRkRlDb0HDNHO0CHPRMDHCRNsOoFMsMkC0DHNRMoCC0sNFRs#VRFsdL.-HR0
RRRRR-RR-RRRRRRRRRRRRNbD0sVFl
#3RRRRRRRR-R-
RRRRR-RR-RRRRRRRR2RLRVACFRsC0RECV#Hs0NROD0DRFhRzQ)wmv0,RE#CRCRC8PkNDCR#
RRRRR-RR-RRRRRRRRRRRR 51 ,74R 1 7R.2ECNPRR0FLHCRMHH0NxDHC08RFNRPD#kCRRHM0RECsoNMCR
RRRRRR-R-RRRRRRRRRRRRrR4,.(4cc6UdnR.9NRM8rR4,.(4ccdUdgRU9sbC#CHO0P$CD3aRRERC
RRRRR-RR-RRRRRRRRRRRRC#C8NRPD#kCRCNsR8lFHCVH8VRN0RCsCENORDONDFR0RQzhwvm)3R
RRRRRR-R-
RRRRRRRRR--RRRRRRRROa2RERH#s8NMFMlRkClLsCRoMNCs0RFsHb#RFNs0LRDCVRFsdL.-HR0
RRRRR-RR-RRRRRRRRRRRRlOFbCk0sR#,NRM8HE0RNN#RRsbCHRF8F~VR.j3d6*Uc5*4j*24URsVFROCNER
RRRRRR-R-RRRRRRRRRRRR#RC0F#VRCRC8PkNDC
#3RRRRRRRR-R-
RRRRR-RR-RRRRRRRR2R8RswFRVHMFNsl0MHFRRFM#ObC0DsNR#0C0V#RF0sRENCRDsoFHl0E,CRsV
CsRRRRRRRR-R-RRRRRRRRRRFR0RC0ER p'OCk$ssRN0DHOC
3
RRRRVOkM0MHFR)BAaXR5RH:RM R)q2pRR0sCkRsM)p q;R
RRRRRR-R-RsukbCF#:R
RRRRRR-R-RRRRRRRRR0)Ck#sMRLOkCFRsFF0RV
RXRRRRRRRR-1-RbHCONPDRNCDk#R:
RRRRR-RR-RRRRRRRRARB)ja53Rj2=3RjjR
RRRRRR-R-RRRRRRRRR)BAa354j=2RRj43
RRRRRRRRR--RRRRRRRRBaA)53-4j=2RR3-4jR
RRRRRR-R-Rl7FN:HM
RRRRRRRRR--RRRRRRRRXMRHRq) pR
RRRRRR-R-Rs sFOsRFHM80MHF#R:
RRRRR-RR-RRRRRRRRFRhMRC
RRRRR-RR-NR)M:oC
RRRRRRRRR--RRRRRRRRBaA)5RX2Hl#RNC0ElHN0ODND$MRkLMFk8
C8RRRRRRRR-h-RF#0C:R
RRRRRR-R-RRRRRRRRRRN2aRECsOCNEDNLCNRsMRoCFBVRAR)aHN#RbFbsGNHl0$CDRPoHCLMR$R:
RRRRR-RR-RRRRRRRRRRRRRRRR1qA5)BAa25X2=R<R)BAa 5)q]p'Q2t]
R
RRkRVMHO0F"MR*R*"5:XRRRHMQ hat; )R:YRRRHM)p q2CRs0MksRq) pR;
RRRRR-RR-kRus#bFCR:
RRRRR-RR-RRRRRRRRCR)0Mks#RRYbCFIsVRFR=XR=R>RXY**
RRRRRRRRR--1ObCHRNDPkNDC
#:RRRRRRRR-R-RRRRRRXRR*3*jjRR=4;3jR/XR=
RjRRRRRRRR-R-RRRRRRjRR*R*Y=3RjjY;RRj>R3Rj
RRRRR-RR-RRRRRRRR*RX*j43R)=R 5qpXR2;X=R>RRj
RRRRR-RR-RRRRRRRR*R4*=YRRj43
RRRRRRRRR--7NFlH
M:RRRRRRRR-R-RRRRRRXRRRj>R
RRRRRRRRR--RRRRRRRRXRR=jFRVsRRY>3RjjR
RRRRRR-R-RRRRRRRRR<XRRVjRFYsRRj=R3Rj
RRRRR-RR-sR sRFsO8FMHF0HM
#:RRRRRRRR-R-RRRRRR RRsssFRRHVXRR<jMRN8RRY/j=R3Rj
RRRRR-RR-RRRRRRRRsR sRFsHXVRRj=RR8NMR<YR=3RjjR
RRRRRR-R-RM)No
C:RRRRRRRR-R-RRRRRRXRR*R*Y>j=R3Rj
RRRRR-RR-FRh0:C#
RRRRRRRRR--RRRRRRRRNa2REkCRbsbCRkLFMF8RVER0CCRsNNOELRDCsoNMCFRVs*R"*H"R#R
RRRRRR-R-RRRRRRRRRRRRNsbbFlGHND0C$HRoPRCML
$:RRRRRRRR-R-RRRRRRRRRRRRRR*RX*<YR= R)q]p'Q
t]
RRRRMVkOF0HM*R"*5"RXRR:H)MR ;qpR:YRRRHM)p q2CRs0MksRq) pR;
RRRRR-RR-kRus#bFCR:
RRRRR-RR-RRRRRRRRCR)0Mks#RRYbCFIsVRFR=XR=R>RXY**
RRRRRRRRR--1ObCHRNDPkNDC
#:RRRRRRRR-R-RRRRRRXRR*3*jjRR=4;3jR/XR=3RjjR
RRRRRR-R-RRRRRRRRRjj3*R*Y=3RjjY;RRj>R3Rj
RRRRR-RR-RRRRRRRR*RX*j43RX=R;RRX>j=R3Rj
RRRRR-RR-RRRRRRRR3R4jY**R4=R3Rj
RRRRR-RR-FR7lMNH:R
RRRRRR-R-RRRRRRRRR>XRRjj3
RRRRRRRRR--RRRRRRRRXRR=jR3jVRFsYRR>j
3jRRRRRRRR-R-RRRRRRXRRRj<R3VjRFYsRRj=R3Rj
RRRRR-RR-sR sRFsO8FMHF0HM
#:RRRRRRRR-R-RRRRRR RRsssFRRHVXRR<jR3jNRM8Y=R/Rjj3
RRRRRRRRR--RRRRRRRR FsssVRHR=XRRjj3R8NMR<YR=3RjjR
RRRRRR-R-RM)No
C:RRRRRRRR-R-RRRRRRXRR*R*Y>j=R3Rj
RRRRR-RR-FRh0:C#
RRRRRRRRR--RRRRRRRRNa2REkCRbsbCRkLFMF8RVER0CCRsNNOELRDCsoNMCFRVs*R"*H"R#R
RRRRRR-R-RRRRRRRRRRRRNsbbFlGHND0C$HRoPRCML
$:RRRRRRRR-R-RRRRRRRRRRRRRR*RX*<YR= R)q]p'Q
t]
RRRRMVkOF0HMmRptXR5RH:RM R)q2pRR0sCkRsM)p qRR=>"_lsD"Fo;R
RRRRRR-R-RsukbCF#:R
RRRRRR-R-RRRRRRRRR0)Ck#sMR0MNkDsNRoDFN0sHEFlRV
RXRRRRRRRR-1-RbHCONPDRNCDk#R:
RRRRR-RR-RRRRRRRRmRpt354j=2RRjj3
RRRRRRRRR--RRRRRRRRp5mtv]qa_R 2=3R4jR
RRRRRR-R-Rl7FN:HM
RRRRRRRRR--RRRRRRRRXRR>j
3jRRRRRRRR- -RsssFRMOF8HH0F:M#
RRRRRRRRR--RRRRRRRR FsssVRHR<XR=3RjjR
RRRRRR-R-RM)No
C:RRRRRRRR-R-RRRRRRpRRmXt52#RHR0lNENCl0NHODRD$kFMLkCM88R
RRRRRR-R-R0hFC
#:RRRRRRRR-R-RRRRRRNRR2ERaCCRsNNOELRDCsoNMCVRFRtpmRRH#NsbbFlGHND0C$HRoPRCML
$:RRRRRRRR-R-RRRRRRRRRRRRRRmRpt+5j2=R<Rtpm5RX2<p=Rm)t5 'qp]]Qt2R

RVRRk0MOHRFM RXu5:XRRRHM)p qRs2RCs0kM R)q=pR>lR"sG_Cb
";RRRRRRRR-u-RkFsb#
C:RRRRRRRR-R-RRRRRR)RRCs0kMC#R*;*XRCIEsCCRRv=Rq_a] R
RRRRRR-R-RC1bODHNRDPNk:C#
RRRRRRRRR--RRRRRRRR 5Xuj23jR4=R3Rj
RRRRR-RR-RRRRRRRRXR u354j=2RRavq]
_ RRRRRRRR-R-RRRRRR RRX-u5423jRv=Rq_a]4e_m  )_
RRRRRRRRR--RRRRRRRR 5XuX=2RRjj3RsVFR<XR=pR-m)t5 'qp]]Qt2R
RRRRRR-R-Rl7FN:HM
RRRRRRRRR--RRRRRRRRXMRHRq) pkR#O0ERERN0 5XuX<2R= R)q]p'Q
t]RRRRRRRR- -RsssFRMOF8HH0F:M#
RRRRRRRRR--RRRRRRRR FsssVRHR>XRRtpm5q) pQ']t
]2RRRRRRRR-)-RNCMo:R
RRRRRR-R-RRRRRRRRRu X5RX2>j=R3Rj
RRRRR-RR-FRh0:C#
RRRRRRRRR--RRRRRRRRNa2REkCR#DNLCFR8lMNHRRFV RXuHN#RbFbsGNHl0$CDRPoHCLMR$R:
RRRRR-RR-RRRRRRRRRRRRRRRR<XR=mRpt 5)q]p'Q2t]
R
RRkRVMHO0FpMRmRt.5:XRRRHM)p qRs2RCs0kM R)q
p;RRRRRRRR-u-RkFsb#
C:RRRRRRRR-R-RRRRRR)RRCs0kMD#RFsoNHl0ER#LNCRR.FXVR
RRRRRRRRR--1ObCHRNDPkNDC
#:RRRRRRRR-R-RRRRRRpRRm5t.423jRj=R3Rj
RRRRR-RR-RRRRRRRRmRpt..53Rj2=3R4jR
RRRRRR-R-Rl7FN:HM
RRRRRRRRR--RRRRRRRRXRR>j
3jRRRRRRRR- -RsssFRMOF8HH0F:M#
RRRRRRRRR--RRRRRRRR FsssVRHR<XR=3RjjR
RRRRRR-R-RM)No
C:RRRRRRRR-R-RRRRRRpRRm5t.XH2R#NRl0lECNO0HN$DDRLkMF8kMCR8
RRRRR-RR-FRh0:C#
RRRRRRRRR--RRRRRRRRNa2REsCRCENONCLDRMsNoFCRVmRptH.R#bRNbGsFH0lNCRD$oCHPM$RL:R
RRRRRR-R-RRRRRRRRRRRRRRRRp.mt52j+RR<=p.mt5RX2<p=Rm5t.)p q't]Q]
2
RRRRVOkM0MHFRtpmR:5XRRHM)p q;qRA1R :H)MR 2qpR0sCkRsM)p q;R
RRRRRR-R-RsukbCF#:R
RRRRRR-R-RRRRRRRRR0)Ck#sMRoDFN0sHELlRNR#CA q1RRFVXR
RRRRRR-R-RC1bODHNRDPNk:C#
RRRRRRRRR--RRRRRRRRp5mt4,3jR1Aq =2RRjj3
RRRRRRRRR--RRRRRRRRp5mtA q1,qRA1R 2=3R4jR
RRRRRR-R-Rl7FN:HM
RRRRRRRRR--RRRRRRRRXRR>j
3jRRRRRRRR-R-RRRRRRARRqR1 >3RjjR
RRRRRR-R-RRRRRRRRR1Aq =R/Rj43
RRRRRRRRR-- FsssFROM08HH#FM:R
RRRRRR-R-RRRRRRRRRs sFHsRVRRX<j=R3Rj
RRRRR-RR-RRRRRRRRsR sRFsHAVRqR1 <j=R3Rj
RRRRR-RR-RRRRRRRRsR sRFsHAVRqR1 =3R4jR
RRRRRR-R-RM)No
C:RRRRRRRR-R-RRRRRRpRRmXt5,qRA1R 2Hl#RNC0ElHN0ODND$MRkLMFk8
C8RRRRRRRR-h-RF#0C:R
RRRRRR-R-RRRRRRRRRRN2WMECR1Aq RR>4,3jRC0ERNsCOLENDsCRNCMoRRFVpRmtHR#
RRRRR-RR-RRRRRRRRRRRRbNbsHFGlCN0Do$RHMPCR:L$
RRRRRRRRR--RRRRRRRRRRRRRpRRmjt5+A,Rq21 RR<=p5mtXA,Rq21 RR<=p5mt)p q't]Q]A,Rq21 
RRRRRRRRR--RRRRRRRRLW2RERCMjR3j<qRA1< RRj43,ER0CCRsNNOELRDCsoNMCVRFRtpmR
H#RRRRRRRR-R-RRRRRRRRRRbRNbGsFH0lNCRD$oCHPM$RL:R
RRRRRR-R-RRRRRRRRRRRRRRRRp5mt)p q't]Q]A,Rq21 RR<=p5mtXA,Rq21 RR<=p5mtjR+,A q12R

RVRRk0MOHRFMp4mtjXR5RH:RM R)q2pRR0sCkRsM)p q;R
RRRRRR-R-RsukbCF#:R
RRRRRR-R-RRRRRRRRR0)Ck#sMRoDFN0sHELlRNR#C4FjRV
RXRRRRRRRR-1-RbHCONPDRNCDk#R:
RRRRR-RR-RRRRRRRRmRpt54j423jRj=R3Rj
RRRRR-RR-RRRRRRRRmRpt54j4jj32RR=4
3jRRRRRRRR-7-RFHlNMR:
RRRRR-RR-RRRRRRRRRRX>3RjjR
RRRRRR-R-Rs sFOsRFHM80MHF#R:
RRRRR-RR-RRRRRRRRsR sRFsHXVRRR<=j
3jRRRRRRRR-)-RNCMo:R
RRRRRR-R-RRRRRRRRRtpm4Xj52#RHR0lNENCl0NHODRD$kFMLkCM88R
RRRRRR-R-R0hFC
#:RRRRRRRR-R-RRRRRRNRR2ERaCCRsNNOELRDCsoNMCVRFRtpm4HjR#bRNbGsFH0lNCRD$oCHPM$RL:R
RRRRRR-R-RRRRRRRRRRRRRRRRp4mtj+5j2=R<Rtpm4Xj52=R<Rtpm4)j5 'qp]]Qt2R

RVRRk0MOHRFMRh1QRR5X:MRHRq) pRR2skC0s)MR Rqp=">Rl#s_H;M"
RRRRRRRRR--ubksF:#C
RRRRRRRRR--RRRRRRRR)kC0sRM##CHMRRFVXX;RRRHMsHN8N
M#RRRRRRRR-1-RbHCONPDRNCDk#R:
RRRRR-RR-RRRRRRRRQR1h25XRj=R3VjRFXsRR	=R*avq]Q_u,ERICRsC	#RHRRNMQ hat
 )RRRRRRRR-R-RRRRRR1RRQXh52RR=4R3jVRFsXRR=5	c*+*42v]qa__uQm)e _R.,IsECCRR	HN#RMR
RRRRRR-R-RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRQRRhta  R)
RRRRR-RR-RRRRRRRRQR1h25XR-=R4R3jVRFsXRR=5	c*+*d2v]qa__uQm)e _R.,IsECCRR	HN#RMR
RRRRRR-R-RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRQRRhta  R)
RRRRR-RR-FR7lMNH:R
RRRRRR-R-RRRRRRRRRHXRM R)qRp
RRRRR-RR-sR sRFsO8FMHF0HM
#:RRRRRRRR-R-RRRRRRhRRF
MCRRRRRRRR-)-RNCMo:R
RRRRRR-R-RRRRRRRRR1qA5h1Q52X2RR<=4
3jRRRRRRRR-h-RF#0C:R
RRRRRR-R-RRRRRRRRRRN2wRFsDoNsCPsRNCDk#VRFR1qA5,X2Ro8CsCN88ORNONksOH$R#DRNDCFI8
3
RRRRVOkM0MHFRmRB1RR5XRR:H)MR Rqp2CRs0MksRq) p>R=Rs"l_#OF"R;
RRRRR-RR-kRus#bFCR:
RRRRR-RR-RRRRRRRRCR)0Mks#FRO#CHMRRFVXX;RRRHMsHN8N
M#RRRRRRRR-1-RbHCONPDRNCDk#R:
RRRRR-RR-RRRRRRRRmRB125XRj=R3VjRFXsRR5=R.+*	4v2*q_a]umQ_e_ ).I,RECCsRH	R#MRN
RRRRRRRRR--RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRQRRhta  R)
RRRRR-RR-RRRRRRRRmRB125XR4=R3VjRFXsRR5=R.2*	*avq]Q_u,ERICRsC	#RHRRNMQ hat
 )RRRRRRRR-R-RRRRRRBRRmX152RR=-j43RsVFR=XRR*5.	2+4*avq]Q_u,ERICRsC	#RHRRNMQ hat
 )RRRRRRRR-7-RFHlNMR:
RRRRR-RR-RRRRRRRRRRXH)MR 
qpRRRRRRRR- -RsssFRMOF8HH0F:M#
RRRRRRRRR--RRRRRRRRhCFM
RRRRRRRRR--)oNMCR:
RRRRR-RR-RRRRRRRRARq1m5B125X2=R<Rj43
RRRRRRRRR--hCF0#R:
RRRRR-RR-RRRRRRRR2RNRswFRsDNoRCsPkNDCF#RVARq125X,CR8o8sNCN8ROsOkNRO$HN#RDIDFC
83
RRRRMVkOF0HMaRRq5hRXRR:H)MR Rqp2CRs0MksRq) pR;
RRRRR-RR-kRus#bFCR:
RRRRR-RR-RRRRRRRRCR)0Mks#NR0MMoC0VRFRRX;XMRHR8sNH#NM
RRRRRRRRR--1ObCHRNDPkNDC
#:RRRRRRRR-R-RRRRRRaRRqXh52RR=jR3jVRFsXRR=	q*vau]_QI,RECCsRH	R#MRNRaQh )t 
RRRRRRRRR--7NFlH
M:RRRRRRRR-R-RRRRRRXRRRRHM)p qR8NM
RRRRRRRRR--RRRRRRRRX=R/R*5.	2+4*avq]Q_u_ me),_.RCIEs	CRRRH#NQMRhta  R)
RRRRR-RR-sR sRFsO8FMHF0HM
#:RRRRRRRR-R-RRRRRR RRsssFRRHVXRR=5*5.	2+4Rv*Rq_a]umQ_e_ ).R2,IsECCRR	HN#RMR
RRRRRR-R-RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRQRRhta  R)
RRRRR-RR-NR)M:oC
RRRRRRRRR--RRRRRRRRa5qhXH2R#NRl0lECNO0HN$DDRLkMF8kMCR8
RRRRR-RR-FRh0:C#
RRRRRRRRR--RRRRRRRRNw2RFDsRNCsosNRPD#kCRRFVq5A1XR2,8sCoN88CRONOkOsN$#RHRDNDF8IC3R

RVRRk0MOHRFMRBq)1RQh5:XRRRHM)p qRs2RCs0kM R)q
p;RRRRRRRR-u-RkFsb#
C:RRRRRRRR-R-RRRRRR)RRCs0kMH#RMsPC##CRHRMCFXVR
RRRRRRRRR--1ObCHRNDPkNDC
#:RRRRRRRR-R-RRRRRRqRR)QB1h35jj=2RRjj3
RRRRRRRRR--RRRRRRRRq1)BQ4h53Rj2=qRvau]_Qe_m .)_
RRRRRRRRR--RRRRRRRRq1)BQ-h5423jR-=Rv]qa__uQm)e _R.
RRRRR-RR-FR7lMNH:R
RRRRRR-R-RRRRRRRRR1qA5RX2<4=R3Rj
RRRRR-RR-sR sRFsO8FMHF0HM
#:RRRRRRRR-R-RRRRRR RRsssFRRHVq5A1X>2RRj43
RRRRRRRRR--)oNMCR:
RRRRR-RR-RRRRRRRRARq1)5qBh1Q5RX2<v=Rq_a]umQ_e_ ).R
RRRRRR-R-R0hFC
#:RRRRRRRR-R-RRRRRRhRRF
MC
RRRRMVkOF0HMqRR)mBB1XR5RH:RM R)q2pRR0sCkRsM)p q;R
RRRRRR-R-RsukbCF#:R
RRRRRR-R-RRRRRRRRR0)Ck#sMRPHMCCs#R#OFHRMCFXVR
RRRRRRRRR--1ObCHRNDPkNDC
#:RRRRRRRR-R-RRRRRRqRR)mBB1354j=2RRjj3
RRRRRRRRR--RRRRRRRRqB)Bmj153Rj2=qRvau]_Qe_m .)_
RRRRRRRRR--RRRRRRRRqB)Bm-15423jRv=Rq_a]uRQ
RRRRR-RR-FR7lMNH:R
RRRRRR-R-RRRRRRRRR1qA5RX2<4=R3Rj
RRRRR-RR-sR sRFsO8FMHF0HM
#:RRRRRRRR-R-RRRRRR RRsssFRRHVq5A1X>2RRj43
RRRRRRRRR--)oNMCR:
RRRRR-RR-RRRRRRRR3Rjj=R<RBq)B5m1X<2R=qRvau]_QR
RRRRRR-R-R0hFC
#:RRRRRRRR-R-RRRRRRhRRF
MC
RRRRMVkOF0HMqRR)qBahYR5RH:RM R)qRp2skC0s)MR ;qp
RRRRRRRRR--ubksF:#C
RRRRRRRRR--RRRRRRRR)kC0sRM#0RECPkNDCVRFRC0ERoNMDHCRMNRs8MHN#VRFRC0ERHbFMR0
RRRRR-RR-RRRRRRRR354jY,R2I,REEHORRH#HsMRCNO0MDokNOsRF8FsH0MNCR#
RRRRR-RR-bR1CNOHDNRPD#kC:R
RRRRRR-R-RRRRRRRRRBq)a5qhj23jRj=R3Rj
RRRRR-RR-FR7lMNH:R
RRRRRR-R-RRRRRRRRRHYRM R)qRp
RRRRR-RR-sR sRFsO8FMHF0HM
#:RRRRRRRR-R-RRRRRRhRRF
MCRRRRRRRR-)-RNCMo:R
RRRRRR-R-RRRRRRRRR1qA5Bq)a5qhYR22<v=Rq_a]umQ_e_ ).R
RRRRRR-R-R0hFC
#:RRRRRRRR-R-RRRRRRhRRF
MC
RRRRMVkOF0HMqRR)qBahYR5RH:RM R)qRp;XRR:H)MR 2qpR0sCkRsM)p q;R
RRRRRR-R-RsukbCF#:R
RRRRRR-R-RRRRRRRRR0)Ck#sMRC0ERHbsMbOHNPDRNCDkRRFV0RECNDMoCMRHR8sNH#NMR
FVRRRRRRRR-R-RRRRRR0RREbCRF0HMR,5XR,Y2RHIEOHER#MRHROsC0oNMksDNRFOFsM8HN#0C
RRRRRRRRR--1ObCHRNDPkNDC
#:RRRRRRRR-R-RRRRRRqRR)qBah35jjX,R2RR=jR3jHXVRRj>R3Rj
RRRRR-RR-RRRRRRRR)RqBhaq5jj3,2RXRv=Rq_a]uHQRVRRX<3RjjR
RRRRRR-R-RRRRRRRRRBq)a5qhYj,R3Rj2=qRvau]_Qe_m .)_RRHVYRR>j
3jRRRRRRRR-R-RRRRRRqRR)qBah,5YRjj32RR=-avq]Q_u_ me)R_.HYVRRj<R3Rj
RRRRR-RR-FR7lMNH:R
RRRRRR-R-RRRRRRRRRHYRM R)qRp
RRRRR-RR-RRRRRRRRRRXH)MR ,qpR/XR=3RjjERICYMRRj=R3Rj
RRRRR-RR-sR sRFsO8FMHF0HM
#:RRRRRRRR-R-RRRRRR RRsssFRRHVXRR=jR3jNRM8YRR=j
3jRRRRRRRR-)-RNCMo:R
RRRRRR-R-RRRRRRRRRq-vau]_QRR<qa)BqYh5,RX2<v=Rq_a]uRQ
RRRRR-RR-FRh0:C#
RRRRRRRRR--RRRRRRRRhCFM
R
RRkRVMHO0F1MRQRh]5:XRRRHM)p q2CRs0MksRq) pR;
RRRRR-RR-kRus#bFCR:
RRRRR-RR-RRRRRRRRCR)0Mks#$REbLCsFODHRM#HCVRFRRX
RRRRR-RR-bR1CNOHDNRPD#kC:R
RRRRRR-R-RRRRRRRRRh1Q]35jj=2RRjj3
RRRRRRRRR--7NFlH
M:RRRRRRRR-R-RRRRRRXRRRRHM)p q
RRRRRRRRR-- FsssFROM08HH#FM:R
RRRRRR-R-RRRRRRRRRMhFCR
RRRRRR-R-RM)No
C:RRRRRRRR-R-RRRRRR1RRQ5h]XH2R#NRl0lECNO0HN$DDRLkMF8kMCR8
RRRRR-RR-FRh0:C#
RRRRRRRRR--RRRRRRRRNa2REkCR#DNLCFR8lMNHRRFV1]QhRRH#NsbbFlGHND0C$HRoPRCML
$:RRRRRRRR-R-RRRRRRRRRRRRRRARq125XRR<=p5mt)p q't]Q]
2

RRRRMVkOF0HMmRB15]RXRR:H)MR 2qpR0sCkRsM)p q;R
RRRRRR-R-RsukbCF#:R
RRRRRR-R-RRRRRRRRR0)Ck#sMRbE$CFsLDRHOOHF#MFCRV
RXRRRRRRRR-1-RbHCONPDRNCDk#R:
RRRRR-RR-RRRRRRRRmRB1j]53Rj2=3R4jR
RRRRRR-R-Rl7FN:HM
RRRRRRRRR--RRRRRRRRXMRHRq) pR
RRRRRR-R-Rs sFOsRFHM80MHF#R:
RRRRR-RR-RRRRRRRRFRhMRC
RRRRR-RR-NR)M:oC
RRRRRRRRR--RRRRRRRRB]m15RX2>4=R3Rj
RRRRR-RR-FRh0:C#
RRRRRRRRR--RRRRRRRRNa2REkCR#DNLCFR8lMNHRRFVB]m1RRH#NsbbFlGHND0C$HRoPRCML
$:RRRRRRRR-R-RRRRRRRRRRRRRRARq125XRR<=p5mt)p q't]Q]
2
RRRRVOkM0MHFRhaq]XR5RH:RM R)qRp2skC0s)MR ;qp
RRRRRRRRR--ubksF:#C
RRRRRRRRR--RRRRRRRR)kC0sRM#EC$bsDLFH0ORNCMoMF0RV
RXRRRRRRRR-1-RbHCONPDRNCDk#R:
RRRRR-RR-RRRRRRRRqRahj]53Rj2=3RjjR
RRRRRR-R-Rl7FN:HM
RRRRRRRRR--RRRRRRRRXMRHRq) pR
RRRRRR-R-Rs sFOsRFHM80MHF#R:
RRRRR-RR-RRRRRRRRFRhMRC
RRRRR-RR-NR)M:oC
RRRRRRRRR--RRRRRRRRq5A1a]qh52X2RR<=4
3jRRRRRRRR-h-RF#0C:R
RRRRRR-R-RRRRRRRRRMhFCR

RVRRk0MOHRFMq1)BQRh]5:XRRRHM)p q2CRs0MksRq) pR;
RRRRR-RR-kRus#bFCR:
RRRRR-RR-RRRRRRRRCR)0Mks#MRHP#CsC$REbLCsFODHRM#HCVRFRRX
RRRRR-RR-bR1CNOHDNRPD#kC:R
RRRRRR-R-RRRRRRRRRBq)1]Qh5jj32RR=j
3jRRRRRRRR-7-RFHlNMR:
RRRRR-RR-RRRRRRRRRRXH)MR 
qpRRRRRRRR- -RsssFRMOF8HH0F:M#
RRRRRRRRR--RRRRRRRRhCFM
RRRRRRRRR--)oNMCR:
RRRRR-RR-RRRRRRRR)RqBh1Q]25XRRH#lEN0C0lNHDONDk$RMkLFM88C
RRRRRRRRR--hCF0#R:
RRRRR-RR-RRRRRRRR2RNRCaERNsCOLENDsCRNCMoRRFVq1)BQRh]HN#RbFbsGNHl0$CDRPoHCLMR$R:
RRRRR-RR-RRRRRRRRRRRRRRRR1qA5Bq)1]Qh52X2RR<=p5mt)p q't]Q]
2
RRRRVOkM0MHFRBq)B]m1RR5X:MRHRq) ps2RCs0kM R)q
p;RRRRRRRR-u-RkFsb#
C:RRRRRRRR-R-RRRRRR)RRCs0kMH#RMsPC#ECR$sbCLHFDOFRO#CHMRRFVXR
RRRRRR-R-RC1bODHNRDPNk:C#
RRRRRRRRR--RRRRRRRRqB)Bm51]423jRj=R3Rj
RRRRR-RR-FR7lMNH:R
RRRRRR-R-RRRRRRRRR>XR=3R4jR
RRRRRR-R-Rs sFOsRFHM80MHF#R:
RRRRR-RR-RRRRRRRRsR sRFsHXVRR4<R3Rj
RRRRR-RR-NR)M:oC
RRRRRRRRR--RRRRRRRRqB)Bm51]X>2R=3RjjR
RRRRRR-R-R0hFC
#:RRRRRRRR-R-RRRRRRNRR2ERaCbRkbRCsLMFk8VRFRC0ERNsCOLENDsCRNCMoRRFVqB)BmR1]HR#
RRRRR-RR-RRRRRRRRRRRRbNbsHFGlCN0Do$RHMPCR:L$RqRR)mBB1X]52=R<Rtpm5q) pQ']t
]2
RRRRMVkOF0HM)RqBhaq]XR5RH:RM R)qRp2skC0s)MR ;qp
RRRRRRRRR--ubksF:#C
RRRRRRRRR--RRRRRRRR)kC0sRM#HCMPsR#CEC$bsDLFH0ORNCMoMF0RV
RXRRRRRRRR-1-RbHCONPDRNCDk#R:
RRRRR-RR-RRRRRRRR)RqBhaq]35jj=2RRjj3
RRRRRRRRR--7NFlH
M:RRRRRRRR-R-RRRRRRqRRAX152RR<4
3jRRRRRRRR- -RsssFRMOF8HH0F:M#
RRRRRRRRR--RRRRRRRR FsssVRHR1qA5RX2>4=R3Rj
RRRRR-RR-NR)M:oC
RRRRRRRRR--RRRRRRRRqa)Bq5h]XH2R#NRl0lECNO0HN$DDRLkMF8kMCR8
RRRRR-RR-FRh0:C#
RRRRRRRRR--RRRRRRRRNa2REsCRCENONCLDRMsNoFCRV)RqBhaq]#RHRbNbsHFGlCN0Do$RHMPCR:L$
RRRRRRRRR--RRRRRRRRRRRRRqRRAq15)qBahX]52<2RRtpm5q) pQ']t
]2
kSVMHO0FPMR_sOF8_HOlCF8_0sFNF0HMj5X:CRsNRD;Y:jRRNsCDZ;RjRR:sDCN;S
SMRR:MkN0s;NDR0sCRM:RNs0kNRD2skC0s)MR Rqp=">RO8FsHlO_F_8CsNF00MHF"
;
CRM8Ravq] _)q
p;
ObN	CNoR8LF$qRva)]_ RqpH
#
RRRR-R-
R-RR-FRpORNDB#FM00NM#FRVs#RzCMRHRC0EROuN	CNoR8AF$MRmDR$
R-RR-R
RRFROMN#0MR0Rv]qa_u _.RR:Rq) p=R:Rd(3U6gj_gnjUdg_jjn6;RRR-C-R*
*.RRRRO#FM00NMRqRvXm_Bz:haRaQh )t RR:=4;6jRR--vHNGlRklOMFk0FRVskRMlsLCRRFV0CsH#R
RRFROMN#0MR0Rv]qa_t Q]ua_QRR:)p qRR:=.463dc.(_.4.U4(_U6dc_(gj(4j_4R6;-*-UbRH
RORRF0M#NRM0RXvq_ Qa)R:RQ hatR ):.=R(R;R-v-RNlGHkblRsHCO#MHFROVN0RFsVRFsO8FsHRO
RORRF0M#NRM0Ravq]__ uR4j:)RR Rqp:.=R.nj.36cn(cg_U(jn_;4(RR--C4**jR
RRFROMN#0MR0Ri:BRRq) p=R:Rjn3(..6gjd6jUUU4Cc.-;j4RR--B#FM00NMRsVFRsOF8
HORRRRO#FM00NMRqRA1  _uR1:)p qRR:=jj3jj;j4R-R-ROwN0RFsVRFsOPFMCCsoMROCO0sHCNsH
R
RR-R-
RRRRR--pNFOD$Rab7CRCNODsHN0FRM#VRFsB8FsHmORbNCs0MHF#R
RR-R-
RRRRb0$CmRB)B7Q_7vm Y_auH R#)R5maaqQ,mhRBe aQm)h;t2
RRRRb0$C R)qep_ mBa)#RHRsNsN5$Rhzqa)RqpsoNMC>R<2VRFRq) pR;
R0RR$RbChzqa)_qpea BmH)R#sRNsRN$5ahqzp)qRMsNo<CR>F2RVqRhaqz)pR;
R#RRk$L0b)CR _qpq_)).#RHRq) p _eB)amRR5j04FR2R;
R#RRk$L0b)CR _qpq_))d#RHRq) p _eB)amRR5j0.FR2R;
R#RRk$L0b)CR _qpea Bmh)_RRH#)p q_Be aRm)50jRFqRvXa_Q ;)2
RRRRL#k0C$bRqTz7h)qa#RHRaQh )t RMsNojCRRR0Fd
;
RRRR-R-
R-RR-kRqGHHDNRs$wOkM0MHF#FRVsFRBsO8HRoqDF0sHE
l#RRRR-R-
RVRRk0MOHRFMu mW)w_m_1._  )Q17R5RH:RMqRhaqz)p _eB)am;hRQQqaQpq_epRz :MRHRq) pR;
RRRRRRRRRRRRRhRRz vA)w_m_peqzR 1:MRHRahqzp)q2CRs0MksRq) p _eB)amR
H#RRRRRRRR-7-RCs#OHHb0F
M:RRRRRRRR-R-RRRRRRCR)0Mks#FRbIRCsF0VRIVFRFNsRROPC0RFsFPVRNCDk#R
RRRRRR-R-R0hFC
#:RRRRRRRR-R-RRRRRRFRhMRC
RRRRR-RR-R
RRRRRRNRPsLHNDeCRR):R _qpea Bm5)RjFR0RvhzA_ )mew_q pz1
2;RRRRRRRRPHNsNCLDRva uRR:)p qRR:=QahQQ_qpezqp R;
RRRRRPRRNNsHLRDCwtpqRA:Rm mpq:hR=)Raz
 ;RRRRLHCoMR
RRRRRRRRRRRRRVRFsQMRHR0jRFzRhv)A __mwezqp D1RF
FbRRRRRRRRRRRRRRRRRQe52=R:Rva uR;
RRRRRRRRRRRRRRRRVRFsuMRHR)7'q htRFDFbR
RRRRRRRRRRRRRRRRRRRRRRRRRRVRHR=QRRu752ER0CRM
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRwRRpRqt:w=Rq p1;R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRGRCH
0;RRRRRRRRRRRRRRRRRRRRRRRRRRRRCRM8H
V;RRRRRRRRRRRRRRRRR8CMRFDFbR;
RRRRRRRRRRRRRRRRHwVRpRqt0MEC
RRRRRRRRRRRRRRRRRRRRRRRRRRRRva u=R:Rva u3/.jR;
RRRRRRRRRRRRRRRRCRM8H
V;RRRRRRRRRRRRRRRRRqwpt=R:Rza) R;
RRRRRRRRRRRRR8CMRFDFbR;
RRRRRRRRRRRRR0sCkRsMeR;
RCRRMu8Rm)W __mw. _1)1Q ;


RRRRO#FM00NMRmaW__qavzQh1RR:)p q_Be aRm):u=Rm)W __mw. _1)1Q 5R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRahqzp)q_Be a'm)5j4j,jRg23,4jR,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRXvq_ Qa)
2;
RRRRMOF#M0N0uR 1mQphRR:)p q_Be a_m)h=R:RR5
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR(RR3dU6gnU4d(dgc.cU(jC-4R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRcRR3nndcj(ngjjjUjjnnjC-4R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR.RR3gcc(nUndn4.U4ncdjC-4R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR4RR3d.c6gcgcn6c(cn4cjC-4R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRnRR34.cUgUjggg666(d4jC-.R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRdRR3d4.gdUdc.djn(U.(jC-.R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR4RR3.6ndU(.nc.j(dnUjjC-.R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR(RR3.U4djc4njj44444njC-dR,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRdRR3ngj.4djdn4gn4g((jC-dR,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR4RR3dg646..4(ncUUU4gjC-dR,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRgRR36(nnU.4gg66dd4g(jC-cR,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRcRR3.UUU44.4c4gU.gUgjC-cR,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR.RR34ccc.jnjg4cd(n46jC-cR,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR4RR3j..(4jd4dUgn.(j4jC-cR,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRnRR3d4j6n464.(cjnU(UjC-6R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRdRR34j6(U6(4646.gnjdjC-6R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR4RR366.Ug(Ujdn44n6(jjC-6R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR(RR3gn.d6gcdj444ggngjC-nR,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRdRR3cU4n.g(nj6nnncgjjC-nR,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR4RR3(gjdncUd4.Uj(4UjjC-nR,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRgRR3n6d(4cdn6cjgUnjjjC-(R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRcRR3U(nd6(4Ud.jj(UUnjC-(R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR.RR3cdU4(U6g44j6j6U4jC-(R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR4RR3.4gjUg.gj66(nUj(jC-(R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR6RR3jgnccnc(d(6g6j6djC-UR,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR.RR3jgU..d.dnU(gj6ddjC-UR,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR4RR3jcg444n4Ugdc6(ncjC-UR,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR(RR3jc666Ujg.ngdUU.4jC-gR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR
2;
RRRRMVkOF0HMmRB)B7QRX5RjRR:H)MR ;qp
RRRRRRRRRRRRRRRRRRRRYRRjRR:H)MR ;qp
RRRRRRRRRRRRRRRRRRRRZRRjRR:H)MR ;qp
RRRRRRRRRRRRRRRRRRRRhRRRH:RMqRhaqz)pR;RRRRRRRRRRRRRR-RR-uRRsHCO#MHFROVN0
FsRRRRRRRRRRRRB7m)QvB_mR7 :MRHR)Bm7_QBv m7_uaY RRRRRRRR-R-RFR)0HN0F5MRZ>R-R
j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RsRFROPC0HFsM5oRY>R-R
j2RRRRRRRRRRRRRRRRRRRR2CRs0MksRq) p)_q)R_dHR#
RRRRR-RR-CR7#HOsbF0HMR:
RRRRR-RR-RRRRRRRRlBFbCk0RsOF8RHOPkNDCR#
RRRRR-RR-FRh0:C#
RRRRRRRRR--RRRRRRRRhCFM
RRRRRRRRRRRRNRPsLHNDXCRR):R Rqp:X=RjR;
RRRRRRRRRRRRPHNsNCLDR:YRRq) p=R:R;Yj
RRRRRRRRRRRRNRPsLHNDZCRR):R Rqp:Z=RjR;
RRRRRRRRRRRRPHNsNCLDRaX_ Rvu: R)q
p;RRRRLHCoMR
RRRRRRRHVB7m)QvB_mR7 =mR)aQqam0hRE
CMRRRRRRRRRVRRFisRRRHMjFR0RDhRF
FbRRRRRRRRRRRRRRRRRRRRR_RXau vRR:=XR;
RRRRRRRRRRRRRRRRRRRRRRHV5RRZ>j=R3Rj20MEC
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRX=R:R-XRR*YRRmaW__qavzQh125i;R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRR:YR=RRY+_RXau vRa*RWqm_aQ_vh5z1i
2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRZRRRR:=ZRR- Qu1p5mhi
2;RRRRRRRRRRRRRRRRRRRRRDRC#RC
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRX:X=RRY+RRa*RWqm_aQ_vh5z1i
2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRYRRRR:=YRR-X _av*uRRmaW__qavzQh125i;R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRR:ZR=RRZ+uR 1mQph25i;R
RRRRRRRRRRRRRRRRRRRRRCRM8H
V;RRRRRRRRRRRRCRM8DbFF;R
RRRRRRDRC#RC
RRRRRRRRRVRRFisRRRHMjFR0RDhRF
FbRRRRRRRRRRRRRRRRRRRRX _av:uR=;RX
RRRRRRRRRRRRRRRRRRRRRHV5RRY<3Rjj02RE
CMRRRRRRRRRRRRRRRRRRRRRRRRRRRRRXRRRR:=XRR-YRR*a_Wmqva_Q1hz5;i2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRY=R:R+YRRaX_ Rvu*WRama_q_hvQzi152R;
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRZ:Z=RR -Rup1Qmih52R;
RRRRRRRRRRRRRRRRRCRRD
#CRRRRRRRRRRRRRRRRRRRRRRRRRRRRRXRRRR:=XRR+YRR*a_Wmqva_Q1hz5;i2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRY=R:R-YRRaX_ Rvu*WRama_q_hvQzi152R;
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRZ:Z=RR +Rup1Qmih52R;
RRRRRRRRRRRRRRRRRCRRMH8RVR;
RRRRRRRRRCRRMD8RF;Fb
RRRRRRRR8CMR;HV
RRRRRRRR0sCkRsM)p q_)q)_5d'XY,R,2RZ;R
RRMRC8mRB)B7Q;R

R-RR-R
RR-R-R8AFHRC#VRFstLDFNvDRNC0ElHN0ORNDwOkM0MHF#0R1NRs0]CCs
RRRR
--RRRRVOkM0MHFRt1QhXR5:MRHRq) pRR2skC0s)MR RqpHR#
RRRRR-RR-CR7#HOsbF0HMR:
RRRRR-RR-RRRRRRRRC1CRMVkOF0HMCR8OsDNNF0HMMRHR Q  0R18jR4(.n3-g4gnR
RRRRRR-R-R0hFC
#:RRRRRRRR-R-RRRRRRFRhMRC
RLRRCMoH
RRRRRRRRRRRHRVR5RRX>3RjjRR2RC0EMR
RRRRRRRRRRRRRRCRs0MksRj43;R
RRRRRRRRRR#CDH5VRR<XRRjj3RR2R0MEC
RRRRRRRRRRRRRRRR0sCkRsM-j43;R
RRRRRRRRRR#CDCR
RRRRRRRRRRRRRRCRs0MksRjj3;R
RRRRRRRRRR8CMR;HV
RRRR8CMRt1Qh
;
RRRRVOkM0MHFRQB pXR5RH:RM R)q2pRR0sCkRsM)p qR
H#RRRRRRRR-7-RCs#OHHb0F
M:RRRRRRRR-R-RRRRRRCR1CkRVMHO0F8MRCNODsHN0FHMRM RQ 1 R048Rj3(n.g-4gRn
RRRRR-RR-FRh0:C#
RRRRRRRRR--RRRRRNRR2FRhRMOFP#CsHRFM0NFRMhRQa  t)$R0bHCR#GRCb0COCR8,#0FRsOkMN
0CRRRRRRRR-R-RRRRRRRRRRMONMRF0FsPCVIDFRsVFRsDNoNCRslokC#M0
RRRRRRRRR--RRRRRLRR2ERaCFR8lMNHRb#kb0FsCL8R$ER0HV#Rk0MOHRFMHX#RRR<=ptq) R
RRRRRR-R-RRRRRRRRO)2RCs0kMX#RRRHVq5A1X>2R=qRp)
t 
RRRRRRRRMOF#M0N0qRp):t Rq) p:RR= R)qQp5hta  ])'Q2t];R
RRRRRRNRPsLHND)CR7):R ;qp
R
RRCRLo
HMRRRRRRRRRRHVq5A1X>2R=qRp)Rt 0MEC
RRRRRRRRRRRRRRRskC0sXMR;R
RRRRRRCRRMH8RV
;
RRRRRRRRRR)7:)=R Rqp5hRQa  t)25X2R;
RRRRRRRRH)VR7RR=XER0CRM
RRRRRRRRRsRRCs0kM7R);R
RRRRRRCRRMH8RV
;
RRRRRRRRRRRRHXVRRj>R30jRE
CMRRRRRRRRRRRRRRRRRRRRRHRRV7R)RR>=XER0CRM
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR0sCkRsM)
7;RRRRRRRRRRRRRRRRRRRRRCRRD
#CRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRCRs0MksRR)7+3R4jR;
RRRRRRRRRRRRRRRRRRRRRMRC8VRH;R
RRRRRRRRRRDRC#RHVR=XRRjj3RER0CRM
RRRRRRRRRRRRRsRRCs0kM3RjjR;
RRRRRRRRRCRRD
#CRRRRRRRRRRRRRRRRRRRRRHRRV7R)RR<=XER0CRM
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR0sCkRsM)+7RRj43;R
RRRRRRRRRRRRRRRRRRRRRR#CDCR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRskC0s)MR7R;
RRRRRRRRRRRRRRRRRRRRRMRC8VRH;R
RRRRRRRRRRMRC8VRH;R
RRMRC8 RBQ
p;
RRRRMVkOF0HMpRwmRm)5:XRRRHM)p qRs2RCs0kM R)qHpR#R
RRRRRR-R-R#7CObsH0MHF:R
RRRRRR-R-RRRRRRRR1RCCVOkM0MHFRO8CDNNs0MHFRRHMQ   R810R(4jn-3.4ngg
RRRRRRRRR--hCF0#R:
RRRRR-RR-RRRRRRRRRN2hOFRFCMPsF#HMFR0RRNMQ hatR )0C$bRRH#CCGbO80C,FR#Rk0sM0ONCR
RRRRRR-R-RRRRRRRRRORRNFMM0PRFCDsVFVIRFDsRNCsoRoNskMlC0R#
RRRRR-RR-RRRRRRRRRL2aREC8NFlH#MRkFbbs80CRRL$0#EHRMVkOF0HM#RHR1qA5RX2<p=Rq )t
RRRRRRRRR--RRRRRORR2CR)0Mks#RRXHqVRAX152=R>R)pqt
 
RRRRRRRRO#FM00NMR)pqtR :)p qR=R:Rq) ph5Qa  t)Q']t;]2
RRRRRRRRsPNHDNLC7R): R)q
p;
RRRRoLCHRM
RRRRRHRRVARq1X5RR>2R=qRp)Rt 0MEC
RRRRRRRRRRRRRRRRRRRR0sCkRsMXR;
RRRRRCRRMH8RV
;
RRRRRRRR):7R= R)q5pRRaQh )t 52X2;R
RRRRRRVRHRR)7=RRX0MEC
RRRRRRRRRRRRRRRR0sCkRsM)
7;RRRRRRRRCRM8H
V;
RRRRRRRRRHVXRR>jR3j0MEC
RRRRRRRRRRRRRRRRRRRRHRRV7R)RR<=XER0CRM
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR0sCkRsM)
7;RRRRRRRRRRRRRRRRRRRRRCRRD
#CRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRCRs0MksRR)7-3R4jR;
RRRRRRRRRRRRRRRRRRRRRMRC8VRH;R
RRRRRRDRC#RHVR=XRRjj3RER0CRM
RRRRRRRRRRRRRsRRCs0kM3RjjR;
RRRRRCRRD
#CRRRRRRRRRRRRRRRRRHRRV7R)RR>=XER0CRM
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR0sCkRsM)-7RRj43;R
RRRRRRRRRRRRRRRRRR#CDCR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRskC0s)MR7R;
RRRRRRRRRRRRRRRRRMRC8VRH;R
RRRRRRMRC8VRH;R
RRMRC8pRwm;m)
R
RRkRVMHO0F)MRm7zhRR5X:MRHRq) pRR2skC0s)MR RqpHR#
RRRRR-RR-CR7#HOsbF0HMR:
RRRRR-RR-RRRRRRRRC1CRMVkOF0HMCR8OsDNNF0HMMRHR Q  0R18jR4(.n3-g4gnR
RRRRRR-R-R0hFC
#:RRRRRRRR-R-RRRRRRNRR2CR)0Mks#3RjjVRHR=XRRjj3
RRRRRRRRR--RRRRRRRRL)2RCs0kMw#Rp)mm5+XRR6j32VRHR>XRRRj
RRRRR-RR-RRRRRRRR2ROR0)Ck#sMRQB pR5X-3Rj6H2RVRRX<
Rj
RRRRoLCHRM
RRRRRRRRRVRHRRRX>3Rjj0RRE
CMRRRRRRRRRRRRRRRRskC0swMRp)mm5+XRR6j32R;
RRRRRRRRRDRC#RHVR<XRRjj3RER0CRM
RRRRRRRRRRRRRsRRCs0kM RBQRp5XRR-j236;R
RRRRRRRRRR#CDCR
RRRRRRRRRRRRRRCRs0MksRjj3;R
RRRRRRRRRR8CMR;HV
RRRR8CMRz)mh
7;
RRRRMVkOF0HM)RazRhB5:XRRRHM)p qRs2RCs0kM R)qHpR#R
RRRRRR-R-R#7CObsH0MHF:R
RRRRRR-R-RRRRRRRR1RCCVOkM0MHFRO8CDNNs0MHFRRHMQ   R810R(4jn-3.4ngg
RRRRRRRRR--hCF0#R:
RRRRR-RR-RRRRRRRR2RNR0)Ck#sMRjj3RRHVXRR=j
3jRRRRRRRR-R-RRRRRRLRR2CR)0Mks#pRwm5m)XH2RVRRX>
RjRRRRRRRR-R-RRRRRRORR2CR)0Mks# RBQXp52VRHR<XRR
j
RRRRLHCoMR
RRRRRRRRRRRHVR>XRRjj3RER0CRM
RRRRRRRRRRRRRsRRCs0kMpRwm5m)X
2;RRRRRRRRRCRRDV#HRRRX<3Rjj0RRE
CMRRRRRRRRRRRRRRRRskC0sBMR 5QpR;X2
RRRRRRRRRRRCCD#
RRRRRRRRRRRRRRRR0sCkRsMj;3j
RRRRRRRRRRRCRM8H
V;RRRRCRM8ah)zB
;

R

RVRRk0MOHRFM"7vm"XR5,:RYRRHM)p qRs2RCs0kM R)qHpR#R
RRRRRR-R-R#7CObsH0MHF:R
RRRRRR-R-RRRRRRRR1RCCVOkM0MHFRO8CDNNs0MHFRRHMQ   R810R(4jn-3.4ngg
RRRRRRRRR--hCF0#R:
RRRRR-RR-RRRRRRRRRN2)kC0sRM#jR3jFCMRsssF
R
RRRRRRNRPsLHNDXCRhq ta QeRA:Rm mpq:hR=RRX<3RjjR;
RRRRRPRRNNsHLRDCYth qeaQ RR:Apmm Rqh:Y=RRj<R3
j;RRRRRRRRPHNsNCLDRpeqz: RRq) pR;
RLRRCMoH
RRRRRRRRR--BOEC	NRPDHH80F$RVMRHbRk0Nksol0CM#R
RRRRRRRRRRVRHRR5Y=3Rjj02RE
CMRRRRRRRRRRRRRRRRR#N#CRs0w1qp R
RRRRRRRRRRRRRRRRRRRRRRCRsb0FsRm"v7,5XRjj32#RHR8kMCMVHC
8"RRRRRRRRRRRRRRRRRRRRRRRR#CCPs$H0R) )m
);RRRRRRRRRRRRRRRRR0sCkRsMj;3j
RRRRRRRRRRRRCRRMH8RV
;
RRRRRRRR-B-RFklb0PCRNCDk
RRRRRRRRRHV5hRX atqQRe 2ER0CRM
RRRRRRRRRRRRRHRRVRR5Yth qeaQ RR20MEC
RRRRRRRRRRRRRRRRRRRRRRRRpeqz: R=RRX+wR5p)mm51qA5/X2q5A1Y222*1qA5;Y2
RRRRRRRRRRRRRRRR#CDCR
RRRRRRRRRRRRRRRRRRRRRRqRepRz :X=RR5+RBp Q51qA5/X2q5A1Y222*1qA5;Y2
RRRRRRRRRRRRRRRR8CMR;HV
RRRRRRRR#CDCR
RRRRRRRRRRRRRRVRHRY5Rhq ta QeR02RE
CMRRRRRRRRRRRRRRRRRRRRRRRRezqp =R:R-XRR 5BQqp5AX152A/q125Y2q2*AY152R;
RRRRRRRRRRRRRCRRD
#CRRRRRRRRRRRRRRRRRRRRRRRRezqp =R:R-XRRp5wm5m)q5A1Xq2/AY152*22q5A1Y
2;RRRRRRRRRRRRRRRRCRM8H
V;RRRRRRRRCRM8H
V;
RRRRRRRR0sCkRsMezqp R;
RCRRM"8Rv"m7;


RRRRVOkM0MHFRq) pXvqR,5XR:YRRRHM)p qRs2RCs0kM R)qHpR#R
RRRRRR-R-R#7CObsH0MHF:R
RRRRRR-R-RRRRRRRR1RCCVOkM0MHFRO8CDNNs0MHFRRHMQ   R810R(4jn-3.4ngg
RRRRRRRRR--hCF0#R:
RRRRR-RR-RRRRRRRRRN2)p qv5qXX2,YRX=RRCIEMRRX=
RYRRRRRRRR-R-
RLRRCMoH
RRRRRRRRRHVX=R>R0YRE
CMRRRRRRRRRsRRCs0kM;RX
RRRRRRRR#CDCR
RRRRRRRRRR0sCkRsMYR;
RRRRRCRRMH8RVR;
RCRRM)8R vqpq
X;
RRRRMVkOF0HM R)qQpvhXR5,RRY:MRHRq) pRR2skC0s)MR RqpHR#
RRRRR-RR-CR7#HOsbF0HMR:
RRRRR-RR-RRRRRRRRC1CRMVkOF0HMCR8OsDNNF0HMMRHR Q  0R18jR4(.n3-g4gnR
RRRRRR-R-R0hFC
#:RRRRRRRR-R-RRRRRR2RNRq) phvQ5YX,2RR=XERICXMRRY=R
RRRRRRRR
--RRRRLHCoMR
RRRRRRVRHR<XR=RRY0MEC
RRRRRRRRRRRskC0sXMR;R
RRRRRRDRC#RC
RRRRRRRRRCRs0MksR
Y;RRRRRRRRCRM8H
V;RRRRCRM8)p qv;Qh
R

RbRRsCFO8CksRQzhwvm)5sPNHDNLC R1 ,7417  .M:HFRk0uQm1a Qe;sPNHDNLC:RXFRk0)p q2R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRHRR#R
RRRRRR-R-R#7CObsH0MHF:R
RRRRRR-R-RRRRRRRR1RCCVOkM0MHFRO8CDNNs0MHFRRHMQ   R810R(4jn-3.4ngg
RRRRRRRRR--hCF0#R:
RRRRR-RR-RRRRRRRRRN2)kC0sRM#jR3jFCMRsssF
RRRRRRRR
--RRRRRRRRPHNsNCLDRRZ,iQ:Rhta  
);RRRRRRRRPHNsNCLDR a1 R74:hRQa  t)=R:RaQh )t ' 51 274;R
RRRRRRNRPsLHNDaCR17  .RR:Q hatR ):Q=Rhta  5)'17  .
2;RRRRLHCoMR
RRRRRR-R-RCBEOP	RN8DHHR0$FNVRslokC#M0
RRRRRRRRRHV17  4RR>.(4cc6Udn0.RE
CMRRRRRRRRRRRRRRRRNC##sw0Rq p1
RRRRRRRRRRRRRRRRRRRRRRRRbsCFRs0" 1 7>4RRc.4(dcU6Rn.HzMRhmQw)
v"RRRRRRRRRRRRRRRRRRRRRRRR#CCPs$H0R) )m
);RRRRRRRRRRRRRRRRX=R:Rjj3;R
RRRRRRRRRRRRRRCRs0Mks;R
RRRRRRMRC8VRH;R

RRRRRHRRV R1 R7.>4R.cU(cdUdgRC0EMR
RRRRRRRRRRRRRR#RN#0CsRpwq1R 
RRRRRRRRRRRRRRRRRRRRRsRRCsbF01R" . 7R.>R4cc(UgddUMRHRQzhwvm)"R
RRRRRRRRRRRRRRRRRRRRRRCR#PHCs0 $R)))m;R
RRRRRRRRRRRRRRRRX:j=R3
j;RRRRRRRRRRRRRRRRskC0s
M;RRRRRRRRCRM8H
V;
RRRRRRRRR--BbFlkR0CMRCI#8CCRDPNkRC#NRM8bk#C8sF-NFM8lkRMlsLC
RRRRRRRR:iR=1Ra 4 7/n6dn
U;RRRRRRRRa 1 7:4R=jRcjR4c*aR517  4RR-iRR*6ndnU-2RR*iRR.4.4
4;
RRRRRRRRRHVa 1 7<4RRRjR0MEC
RRRRRRRRRRRRRRRR a1 R74:a=R17  4RR+.(4cc6Udn
d;RRRRRRRRCRM8H
V;
RRRRRRRR:iR=1Ra . 7/(6.(
c;RRRRRRRRa 1 7:.R=jRcnRg.*aR517  .RR-iRR*6(.(c-2RR*iRRgd(4
;
RRRRRRRRHaVR17  .RR<j0RRE
CMRRRRRRRRRRRRRRRRa 1 7:.R=1Ra . 7R.+R4cc(UgddgR;
RRRRRCRRMH8RV
;
RRRRRRRRZ=R:R a1 R74-1Ra . 7;R
RRRRRRVRHR<ZRR04RE
CMRRRRRRRRRRRRRRRRZ=R:R+ZRRc.4(dcU6;n.
RRRRRRRR8CMR;HV
R
RRRRRR-R-R0tCR0FkbRk0PkNDCR#
RRRRR1RR 4 7RR:=uQm1a Qe'15a 4 72R;
RRRRR1RR . 7RR:=uQm1a Qe'15a . 72R;
RRRRRXRRRR:=Rq) p25Z*nc364nnd4C-jR;
RCRRMz8RhmQw)
v;
R

RVRRk0MOHRFM1aT)RR5X:MRHRq) pRR2skC0s)MR RqpHR#
RRRRR-RR-CR7#HOsbF0HMR:
RRRRR-RR-RRRRRRRRC1CRMVkOF0HMCR8OsDNNF0HMMRHR Q  0R18jR4(.n3-g4gnR
RRRRRR-R-R0hFC
#:RRRRRRRR-R-RRRRRR2RNRCz##ER0CCRhIM0F-b)NEM#FRbNbsHFGlHN0F
M:RRRRRRRR-R-RRRRRRRRRR5RwM2+4Rj=R3r6*w25MRG+R/Mw52R9
RRRRR-RR-RRRRRRRRRL2)kC0sRM#jR3jFCMRsssF
RRRRRRRR
--
RRRRRRRRMOF#M0N0uR 1RR:)p qRR:=A q1_1 u*1Aq u_ 1-;R-FRBMsPCoOCMCNRVOs0F
R
RRRRRRNRPsLHNDQCRhqQep):R ;qp
RRRRRRRRsPNHDNLCpRm7peqR):R Rqp;R
RRRRRRNRPsLHNDhCR qWepRR:)p qRR;
RRRRRPRRNNsHLRDCBhmzaRR:Q hatR ):4=R;R

RLRRCMoH
RRRRRRRRR--BOEC	NRPDHH80F$RVsRNoCklMR0
RRRRRHRRVRR5XRR<jR3j2ER0CRM
RRRRRRRRRRRRRNRR#s#C0qRwp
1 RRRRRRRRRRRRRRRRRRRRRRRRsFCbs"0RXRR<jR3jH1MRT5)aX
2"RRRRRRRRRRRRRRRRRRRRRRRR#CCPs$H0R) )m
);RRRRRRRRRRRRRRRRskC0sjMR3
j;RRRRRRRRCRM8H
V;
RRRRRRRRR--tRC00REC#NJkssCRFRF0VRFs#ObCHRNDOCN##R
RRRRRRVRHR=XRRjj3RC0EMR
RRRRRRRRRRRRRRRRRskC0sjMR3
j;RRRRRRRRCCD#
RRRRRRRRRRRRRRRRRHV5RRX=3R4jRR20MEC
RRRRRRRRRRRRRRRRRRRRRRRR0sCkRsM4;3j
RRRRRRRRRRRRRRRR8CMR;HV
RRRRRRRR8CMR;HV
R
RRRRRR-R-R0tCRC0ERk#JNRsCs0FFRsVFRMoCCDsNR#ONCR#
RRRRRQRRhqQep=R:Ru X5tpm5*X256j32R2;-v-RNC0ElHN0ODND$FROsOsC0kRL0lRHbOsCH
#CRRRRRRRRmep7q:pR=hRQQpeq;R
RRRRRR RhWpeqRR:=5mX/pq7epRR+mep7q*p2j;36
R
RRRRRR-R-RCBEOV	RFRsRsNCD0CHPR8NMR#NLF0DkCsRCsRFsNRM8lRNGOMFk0R
RRRRRRERIHRDCR55RRA5q1h55 qWepmR-pq7eph2/ qWep>2RR1 u2)Rm
RRRRRRRRRRRRRRRRRRR51qA5Wh eRqp-pRm7peq2RR> 2u1Rq2RhR7
RRRRRRRRRRRRRRRRRBR5mazhRv<RqBX_mazh2RR2RFDFbR
RRRRRRRRRRRRRRpRm7peqRR:=he Wq
p;RRRRRRRRRRRRRRRRhe Wq:pR=XR5/7mpeRqp+pRm7peq23*j6R;
RRRRRRRRRRRRRBRRmazhRR:=BhmzaRR+4R;
RRRRRCRRMD8RF;Fb
RRRRRRRR0sCkRsMhe Wq
p;RRRRCRM81aT);R

RVRRk0MOHRFMBaA)RR5X:MRHRq) pRR2skC0s)MR RqpHR#
RRRRR-RR-CR7#HOsbF0HMR:
RRRRR-RR-RRRRRRRRC1CRMVkOF0HMCR8OsDNNF0HMMRHR Q  0R18jR4(.n3-g4gnR
RRRRRR-R-R0hFC
#:RRRRRRRR-R-RRRRRR2RNRCz##ER0CCRhIM0F-b)NEM#FRbNbsHFGlHN0F
M:RRRRRRRR-R-RRRRRRRRRR5RwM2+4R5=R42/d**r.w25MRG+R/Mw52.**9R;
RRRRR-RR-R
RRRRRRFROMN#0M 0Ru:1RRq) p=R:R1Aq u_ 1q*A1  _u
1;
RRRRRRRRsPNHDNLChRQQpeq: R)q
p;RRRRRRRRPHNsNCLDRmXpBRqp: R)q:pR=;RX
RRRRRRRRsPNHDNLC RhtQqae: RRmAmph qRR:=XRR<j;3j
RRRRRRRRsPNHDNLCpRm7peqR):R Rqp;R
RRRRRRNRPsLHNDhCR qWepRR:)p qRR;
RRRRRPRRNNsHLRDCBhmzaRR:Q hatR ):4=R;R

RLRRCMoH
R
RRRRRR-R-RlBFbCk0RFsF0FRVsbR#CNOHDNRO#
C#RRRRRRRRHXVRRj=R30jRE
CMRRRRRRRRRRRRRRRRskC0sjMR3
j;RRRRRRRRCHD#VRR5XRR=4R3j2ER0CRM
RRRRRRRRRRRRRsRRCs0kM3R4jR;
RRRRRCRRD
#CRRRRRRRRRRRRRRRRHXVRR-=R4R3j0MEC
RRRRRRRRRRRRRRRRRRRRRRRR0sCkRsM-j43;R
RRRRRRRRRRRRRRMRC8VRH;R
RRRRRRMRC8VRH;R

RRRRR-RR-FRBl0bkCFRsFV0RFosRCsMCNODRN##C
RRRRRRRRRHVhq ta QeRC0EMR
RRRRRRRRRRRRRRpRXmpBqRR:=-
X;RRRRRRRRCRM8H
V;
RRRRRRRRQQheRqp: =RXpu5mXt5pqmBp52/d23j2-;R-NRv0lECNO0HN$DDRsOFs0COR0Lk
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-lRHbOsCH
#CRRRRRRRRmep7q:pR=hRQQpeq;R
RRRRRR RhWpeqRR:=5mXpB/qp57mpe*qpmep7qRp2+3R.jp*m7peq23/dj
;
RRRRRRRR-B-RE	CORsVFRDsCNP0HCMRN8LRN#kFD0CCRsssF#MRN8NRlGFROk
M0RRRRRRRRIDEHCRR555RRq5A15Wh eRqp-7mpe2qp/Wh e2qpR >Ru21RR
m)RRRRRRRRRRRRRRRRR5RRq5A1he Wq-pRR7mpe2qpR >Ru21RRR2Rq
h7RRRRRRRRRRRRRRRRR5RRRzBmh<aRRXvq_zBmh2aRRD2RF
FbRRRRRRRRRRRRRRRRmep7q:pR= RhWpeq;R
RRRRRRRRRRRRRR RhWpeqR5:=XBpmq5p/mep7qmp*pq7ep+2RRj.3*7mpe2qp/jd3;R
RRRRRRRRRRRRRRmRBzRha:B=RmazhR4+R;R
RRRRRRMRC8FRDF
b;
RRRRRRRRRHVhq ta QeRC0EMR
RRRRRRRRRRRRRR RhWpeqRR:=-Wh e;qp
RRRRRRRR8CMR;HV
R
RRRRRRCRs0MksRWh e;qp
RRRR8CMR)BAa
;
RRRRVOkM0MHFR*"*"XR5RH:RMhRQa  t)Y;RRH:RM R)qRp2skC0s)MR RqpHR#
RRRRR-RR-CR7#HOsbF0HMR:
RRRRR-RR-RRRRRRRRC1CRMVkOF0HMCR8OsDNNF0HMMRHR Q  0R18jR4(.n3-g4gnR
RRRRRR-R-R0hFC
#:RRRRRRRR-R-RRRRRR2RNR0)Ck#sMRjj3RRFMCFsssFROM08HH
FM
RRRRoLCHRM
RRRRR-RR-ERBCRO	PHND8$H0RRFVNksol0CM
RRRRRRRRRHV5RR5XRR<j2RRR8NMRY5RRR/=jR3j2RR20MEC
RRRRRRRRRRRRRRRR#N#CRs0w1qp R
RRRRRRRRRRRRRRRRRRRRRRCRsb0FsRR"X<RRjNRM8Y=R/Rjj3RRHMXY**"R
RRRRRRRRRRRRRRRRRRRRRRCR#PHCs0 $R)))m;R
RRRRRRRRRRRRRRCRs0MksRjj3;R
RRRRRRMRC8VRH;R

RRRRRHRRVRR55RRX=RRjRN2RM58RR<YR=3RjjRR22ER0CRM
RRRRRRRRRRRRRNRR#s#C0qRwp
1 RRRRRRRRRRRRRRRRRRRRRRRRsFCbs"0RXRR=jMRN8RRY<j=R3HjRM*RX*
Y"RRRRRRRRRRRRRRRRRRRRRRRR#CCPs$H0R) )m
);RRRRRRRRRRRRRRRRskC0sjMR3
j;RRRRRRRRCRM8H
V;
RRRRRRRRR--tRC0PkNDCFRVsbR#CNOHDNRO#
C#RRRRRRRRH5VRR=XRRRjRNRM8R>YRRjj3R02RE
CMRRRRRRRRRRRRRRRRskC0sjMR3
j;RRRRRRRRCRM8H
V;
RRRRRRRRRHV5RRX=RR42ER0CRM
RRRRRRRRRRRRRsRRCs0kM3R4jR;
RRRRRCRRMH8RV
;
RRRRRRRRH5VRR=YRRjj3R8NMR/XR=RRj2ER0CRM
RRRRRRRRRRRRRsRRCs0kM3R4jR;
RRRRRCRRMH8RV
;
RRRRRRRRH5VRR=YRRj432ER0CRM
RRRRRRRRRRRRRsRRCs0kM)R5 5qpX;22
RRRRRRRR8CMR;HV
R
RRRRRR-R-R0tCRDPNkVCRFosRCsMCNODRN
#CRRRRRRRRskC0s MRX5uRYRR*pRmt5q) p25X2
2;RRRRCRM8""**;R

RVRRk0MOHRFM""**RR5X:MRHRq) pY;RRH:RM R)qRp2skC0s)MR RqpHR#
RRRRR-RR-CR7#HOsbF0HMR:
RRRRR-RR-RRRRRRRRC1CRMVkOF0HMCR8OsDNNF0HMMRHR Q  0R18jR4(.n3-g4gnR
RRRRRR-R-R0hFC
#:RRRRRRRR-R-RRRRRR2RNR0)Ck#sMRjj3RRFMCFsssFROM08HH
FM
RRRRoLCHRM
RRRRR-RR-ERBCRO	PHND8$H0RRFVNksol0CM
RRRRRRRRRHV5RR5XRR<jR3jRN2RM58RR/YR=3RjjRR22ER0CRM
RRRRRRRRRRRRRNRR#s#C0qRwp
1 RRRRRRRRRRRRRRRRRRRRRRRRsFCbs"0RXRR<jR3jNRM8Y=R/Rjj3RRHMXY**"R
RRRRRRRRRRRRRRRRRRRRRRCR#PHCs0 $R)))m;R
RRRRRRRRRRRRRRCRs0MksRjj3;R
RRRRRRMRC8VRH;R

RRRRRHRRVRR55RRX=3Rjj2RRR8NMRY5RRR<=jR3j2RR20MEC
RRRRRRRRRRRRRRRR#N#CRs0w1qp R
RRRRRRRRRRRRRRRRRRRRRRCRsb0FsRR"X=3RjjMRN8RRY<j=R3HjRM*RX*
Y"RRRRRRRRRRRRRRRRRRRRRRRR#CCPs$H0R) )m
);RRRRRRRRRRRRRRRRskC0sjMR3
j;RRRRRRRRCRM8H
V;
RRRRRRRRR--tRC0PkNDCFRVsbR#CNOHDNRO#
C#RRRRRRRRH5VRR=XRRjj3RMRN8YRRRj>R32jRRC0EMR
RRRRRRRRRRRRRRCRs0MksRjj3;R
RRRRRRMRC8VRH;R

RRRRRHRRVRR5XRR=4R3j2ER0CRM
RRRRRRRRRRRRRsRRCs0kM3R4jR;
RRRRRCRRMH8RV
;
RRRRRRRRH5VRR=YRRjj3R8NMR/XR=3RjjRR20MEC
RRRRRRRRRRRRRRRR0sCkRsM4;3j
RRRRRRRR8CMR;HV
R
RRRRRRVRHRY5RR4=R3Rj20MEC
RRRRRRRRRRRRRRRR0sCkRsM5;X2
RRRRRRRR8CMR;HV
R
RRRRRR-R-R0tCRDPNkVCRFosRCsMCNODRN
#CRRRRRRRRskC0s MRX5uRYRR*pRmt52X2;R
RRMRC8*R"*
";
A--zaQpQ1hz R7RRkRVMHO0F MRXRuR5:XRRRHM)p qRs2RCs0kM R)qHpR#-
-ApzQazQh1R 7RRRRR-RR-CR7#HOsbF0HM-:
-QAzphaQz71 RRRRRRRR-R-RRRRRRCR1CkRVMHO0F8MRCNODsHN0FHMRM RQ 1 R048Rj3(n.g-4g-n
-QAzphaQz71 RRRRRRRR-h-RF#0C:-
-ApzQazQh1R 7RRRRR-RR-RRRRRRRRRN2a#EHRMVkOF0HMFROl0bkC0#RECCRGMbFCHM0NkDR#oHMRC0ERDVFDHFIM-o
-QAzphaQz71 RRRRRRRR-R-RRRRRRRRRRs#CH:C#
A--zaQpQ1hz R7RRRRRR-R-RRRRRRRRRRRRRRRRC5GbG=2RR+4RR+GRR*G*.!/.RG+R*/*dd+!RR333R|;RG<|RRj43
A--zaQpQ1hz R7RRRRRR-R-RRRRRRRRRNRRMs8RCO8kCN#RslokCRM0XFR0R	0NC8RNP0NMNRoCFCVRGGb5+R$2=-
-ApzQazQh1R 7RRRRR-RR-RRRRRRRRRRRC5GbGC2*G$b52-
-ApzQazQh1R 7RRRRR-RR--
-ApzQazQh1R 7RRRRR-RR-RRRRRRRRRL2a#EHRbHlDCClM00NHRFMDHHl0X#RRR0FLDCRCR##0MENRtpm5q) pQ']t
]2-z-AQQpah z17RRRRRRRRR--RRRRRRRRRFR0RFNPHF8RPVCsD3FIRCR)0Mks# R)q]p'QRt]IMECRsXRCENOC0#RE
N0-z-AQQpah z17RRRRRRRRR--RRRRRRRRRHRDl
H0-z-AQQpah z17RRRRRRRR
---z-AQQpah z17RRRRRRRRMOF#M0N0uR 1RR:)p qRR:=A q1_1 u*1Aq u_ 1q*A1  _u-1;-sRuC#OHHRFMO0sHCNsH
A--zaQpQ1hz -7
-QAzphaQz71 RRRRRRRRRRRRPHNsNCLDRB) Qmu)B:qpRmAmph qRR:=XRR<j;3j-B-RE	CORo#HMVRFRoNskMlC0-
-ApzQazQh1R 7RRRRRRRRRPRRNNsHLRDCXBpmq:pRRq) p=R:R1qA5;X2RRRRR-RR-#RzCFRb#HH0PPCRNCDk
A--zaQpQ1hz R7RRRRRRRRRRNRPsLHNDmCRpq7ep):R Rqp;-
-ApzQazQh1R 7RRRRRRRRRPRRNNsHLRDCBhmzaQ:Rhta  ;)R
A--zaQpQ1hz R7RRRRRRRRRRNRPsLHNDhCR qWep):R Rqp;-
-ApzQazQh1R 7RRRRRRRRRPRRNNsHLRDCpaq1_)a v):R Rqp;-
-ApzQazQh1R 7RRRRRPRRNNsHLRDCwaqBm:)RRq) p=R:Rj43;-
-ApzQazQh1
 7-z-AQQpah z17RRRRCRLo
HM-z-AQQpah z17RRRRRRRRRRRRR--BbFlkR0CPkNDCFRVsbR#CNOHDNRO#
C#-z-AQQpah z17RRRRRRRRRHVXRR=jR3j0MEC
A--zaQpQ1hz R7RRRRRRRRRRRRRRCRs0MksRj43;-
-ApzQazQh1R 7RRRRRCRRMH8RV-;
-QAzphaQz71 
A--zaQpQ1hz R7RRRRRRVRHRpRXmpBqR4=R3RjR0MEC
A--zaQpQ1hz R7RRRRRRRRRRRRRRVRHRB) Qmu)BRqp0MEC
A--zaQpQ1hz R7RRRRRRRRRRRRRRRRRRRRRRCRs0MksRavq]__4m)e _
 ;-z-AQQpah z17RRRRRRRRRRRRRRRR#CDC-
-ApzQazQh1R 7RRRRRRRRRRRRRRRRRRRRRsRRCs0kMqRva ]_;-
-ApzQazQh1R 7RRRRRRRRRRRRRCRRMH8RV-;
-QAzphaQz71 RRRRRRRRCRM8H
V;-z-AQQpah z17-
-ApzQazQh1R 7RRRRRHRRVXRRpqmBpRR=.R3jRC0EM-
-ApzQazQh1R 7RRRRRRRRRRRRRHRRV R)B)QumpBqRC0EM-
-ApzQazQh1R 7RRRRRRRRRRRRRRRRRRRRRsRRCs0kM3R4jq/va ]__;u.
A--zaQpQ1hz R7RRRRRRRRRRRRRRDRC#-C
-QAzphaQz71 RRRRRRRRRRRRRRRRRRRRRRRRskC0svMRq_a] ._u;-
-ApzQazQh1R 7RRRRRRRRRRRRRCRRMH8RV-;
-QAzphaQz71 RRRRRRRRCRM8H
V;-z-AQQpah z17-
-ApzQazQh1R 7RRRRRHRRVXRRpqmBpRR=4jj3RER0C-M
-QAzphaQz71 RRRRRRRRRRRRRRRRH)VR uBQ)qmBpER0C-M
-QAzphaQz71 RRRRRRRRRRRRRRRRRRRRRRRRskC0s4MR3vj/q_a] 4_uj-;
-QAzphaQz71 RRRRRRRRRRRRRRRRCCD#
A--zaQpQ1hz R7RRRRRRRRRRRRRRRRRRRRRRCRs0MksRavq]__ u;4j
A--zaQpQ1hz R7RRRRRRRRRRRRRRMRC8VRH;-
-ApzQazQh1R 7RRRRRCRRMH8RV-;
-QAzphaQz71 
A--zaQpQ1hz R7RRRRRRVRHRmXpBRqp>mRpt 5)q]p'Q2t]RC0EM-
-ApzQazQh1R 7RRRRRRRRRRRRRHRRV R)B)QumpBqRC0EM-
-ApzQazQh1R 7RRRRRRRRRRRRRRRRRRRRRsRRCs0kM3Rjj-;
-QAzphaQz71 RRRRRRRRRRRRRRRRCCD#
A--zaQpQ1hz R7RRRRRRRRRRRRRRRRRRRRRR#RN#0CsRpwq1- 
-QAzphaQz71 RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRsFCbs"0RXRR>p5mt)p q't]Q]H2RMXR u25X"-
-ApzQazQh1R 7RRRRRRRRRRRRRRRRRRRRRRRRRRRRR#RRCsPCHR0$h ma;-
-ApzQazQh1R 7RRRRRRRRRRRRRRRRRRRRRsRRCs0kM R)q]p'Q;t]
A--zaQpQ1hz R7RRRRRRRRRRRRRRMRC8VRH;-
-ApzQazQh1R 7RRRRRCRRMH8RV-;
-QAzphaQz71 
A--zaQpQ1hz R7RRRRRR-R-R8)CkROCNksol0CMRR0Fq5A1X<2RRj43
A--zaQpQ1hz R7RRRRRRERIHRDCXBpmq>pRR34jjFRDF-b
-QAzphaQz71 RRRRRRRRRRRRRRRRXBpmq:pR=pRXmpBqR4-Rj;3j
A--zaQpQ1hz R7RRRRRRRRRRRRRRqRwB)amRR:=waqBmv)*q_a] 4_uj-;
-QAzphaQz71 RRRRRRRRCRM8DbFF;-
-ApzQazQh1
 7-z-AQQpah z17RRRRRRRRHIEDXCRpqmBpRR>4R3jDbFF
A--zaQpQ1hz R7RRRRRRRRRRRRRRpRXmpBqRR:=XBpmq-pRRj43;-
-ApzQazQh1R 7RRRRRRRRRRRRRwRRqmBa)=R:RBwqa*m)v]qa_
 ;-z-AQQpah z17RRRRRRRR8CMRFDFb-;
-QAzphaQz71 
A--zaQpQ1hz R7RRRRRR-R-RlBFbCk0RDPNkVCRFOsRNR#CjRR<XBpmq<pRR-4
-QAzphaQz71 RRRRRRRRmep7q:pR=3R4j-;
-QAzphaQz71 RRRRRRRRpaq1_)a v=R:RmXpB;qp
A--zaQpQ1hz R7RRRRRR RhWpeq:m=Rpq7epRR+paq1_)a v-;
-QAzphaQz71 RRRRRRRRBhmza=R:R
.;-z-AQQpah z17-
-ApzQazQh1R 7RRRRR-RR-ERBCRO	VRFssNCD0CHPR8NMR#NLF0DkCsRCs#FsR8NMRGlNRkOFM-0
-QAzphaQz71 RRRRRRRRIDEHCRR55qR5A515he Wq-pRR7mpe2qp/Wh e2qpR >RuR12m-)
-QAzphaQz71 RRRRRRRRRRRRRRRRRqR5Ah15 qWepRR-mep7qRp2>uR 122RR7qh
A--zaQpQ1hz R7RRRRRRRRRRRRRRRRR5zBmh<aRRXvq_zBmh2aRRD2RF
Fb-z-AQQpah z17RRRRRRRRRRRRRRRR7mpeRqp:h=R qWep-;
-QAzphaQz71 RRRRRRRRRRRRRRRRpaq1_)a v=R:R1pqa _a)5v*XBpmq/pRR 5)qBp5mazh2;22
A--zaQpQ1hz R7RRRRRRRRRRRRRR RhWpeqRR:=mep7q+pRR1pqa _a)
v;-z-AQQpah z17RRRRRRRRRRRRRRRRzBmh:aR=mRBzRha+;R4
A--zaQpQ1hz R7RRRRRRMRC8FRDF
b;-z-AQQpah z17-
-ApzQazQh1R 7RRRRR-RR-FRBl0bkCHRVMRNDPkNDC#RkHRMoC5GbG2+$RC=RGGb52G*Cb25$
A--zaQpQ1hz R7RRRRRR RhWpeqRR:=he Wqwp*qmBa)-;
-QAzphaQz71 
A--zaQpQ1hz R7RRRRRRVRHRB) Qmu)BRqp0MEC
A--zaQpQ1hz R7RRRRRRRRRRRRRR RhWpeqRR:=4/3jhe Wq
p;-z-AQQpah z17RRRRRRRR8CMR;HV
A--zaQpQ1hz -7
-QAzphaQz71 RRRRRRRRskC0shMR qWep-;
-QAzphaQz71 RRRRR8CMRu X;


RRRR-R-
R-RR-kRqGHHDNRs$wOkM0MHF#FR0RlBFbCk0Rtpm
RRRR
--RRRRVOkM0MHFRmQptXA5:MRHRq) ps2RCs0kMhRQa  t)1RQ
RRRRRRRRR--7OC#s0HbH:FM
RRRRRRRRR--RRRRR)RRCs0kMM#RRO#kEER0N-0R4=R<R1qA5/X2.R^M<
R.RRRRRRRR-h-RF#0C:R
RRRRRR-R-RRRRRRRRhCFM
R
RRRRRRNRPsLHNDhCR:hRQa  t)=R:R
j;RRRRRRRRPHNsNCLDRRY:)p qRR:=q5A1X
2;
RRRRoLCHRM
RRRRRHRRVR5Y=3R4jsRFR=YRRjj32ER0CRM
RRRRRRRRRRRRRsRRCs0kM;Rj
RRRRRRRR8CMR;HV
R
RRRRRRVRH5RRY>3R4j02RE
CMRRRRRRRRRRRRRRRRIDEHCRRY>.=R3DjRF
FbRRRRRRRRRRRRRRRRRRRRRRRRY=R:R.Y/3
j;RRRRRRRRRRRRRRRRRRRRRRRRh=R:R4h+;R
RRRRRRRRRRRRRRMRC8FRDF
b;RRRRRRRRRRRRRRRRskC0shMR;R
RRRRRRMRC8VRH;R

RRRRR-RR-RRm<RRY<
R4RRRRRRRRIDEHCRRY<3R4jFRDFRb
RRRRRRRRRRRRRYRRRR:=Y3*.jR;
RRRRRRRRRRRRRhRRRR:=h4R-;R
RRRRRRMRC8FRDF
b;RRRRRRRRskC0shMR;R
RRMRC8pRQm;tA
R
RRkRVMHO0FpMR7u X5RX:H)MR ;qpRRh:HQMRhta  R)2)z a))hR RqpQR1
RRRRR-RR-CR7#HOsbF0HMR:
RRRRR-RR-RRRRRRRR0)Ck#sMR.X*^RM
RRRRR-RR-FRh0:C#
RRRRRRRRR--RRRRRRRRhCFM
RRRRoLCHRM
RRRRRsRRCs0kM*RX5j.3RR**h
2;RRRRCRM8pX7 u
;
-z-AQQpah z17RRRRMVkOF0HMmRptXR5RH:RM R)q2pRR0sCkRsM)p qR
Q1-z-AQQpah z17RRRRRRRRR--7OC#s0HbH:FM
A--zaQpQ1hz R7RRRRRR-R-RRRRRRRR1RCCVOkM0MHFRO8CDNNs0MHFRRHMQ   R810R(4jn-3.4ngg
A--zaQpQ1hz R7RRRRRR-R-
A--zaQpQ1hz R7RRRRRR-R-R0hFC
#:-z-AQQpah z17RRRRRRRRR--RRRRRNRR2CR)0Mks# R)qpp'mFWRMsRCs
Fs-z-AQQpah z17RRRRRRRR
---z-AQQpah z17RRRRRRRRR--B$FbsEHo0OR52gR4g).RCMoC0F#RVER0CMRzHsPC#$H0RRFVBHNDVMFsH
N3-z-AQQpah z17RRRRRRRRR--qRDDsEHo0s#RCs#CP3C8
A--zaQpQ1hz R7RRRRRR-R-
A--zaQpQ1hz R7RRRRRR-R-R8)CHs#0H0LkHRFMNRM8kR#CH#MRFOksCMRN8HRLM$NsRsVFlR#,IEH0RRFsIEH0F
k0-z-AQQpah z17RRRRRRRRR--lHF8VNHO0MHF,sRNCCRbs0lH0RC8bPsFH88CRN0E0ER0CFRVDIDFHRMoO8FMHF0HM-#
-QAzphaQz71 RRRRRRRR-N-RslCRC
0:-z-AQQpah z17RRRRRRRRR--4)3RC#8H0LsHkF0HMF#RVFR#kCsOR8OFCkRl#s0RCH0NMER0CLRNFRPCO$FbsEHo0-
-ApzQazQh1R 7RRRRR-RR-FRM0CHO,ER0HD#RHR#0FOVRFHM80MHF#MRN8ER0CFRVDIDFHRMo8OH#DlNHC
s3-z-AQQpah z17RRRRRRRRR--.)3RC#8H0LsHkF0HMH#RMHRLM$NsRsVFlkRl#s0RCFbs8CkORC0ERFNLPOCRFsb$H0oE
A--zaQpQ1hz R7RRRRRR-R-R0MFH,OCRH0E#HRD#F0RVFROM08HH#FMR8NMRC0ERDVFDHFIM8oRHD#ONCHlsMRHRC0E
A--zaQpQ1hz R7RRRRRR-R-RO8FkMlC0HN0FNMRMF8/s0RFERCslCN0sDHN#sRbF8PHCI8RHR0E0REC80H#skHL0MHF3-
-ApzQazQh1R 7RRRRR-RR-3RdRDqDRPN8CHs0#oHMR0lNCNsHDl#RCHM0FMMHoCRVNs0kCF#Rs#RkCVRFRH0E#-
-ApzQazQh1R 7RRRRR-RR-FR#VN0IslCRkR#08bH#DRN$0RECVDFDFMIHoORN	IMFDoC8CMlC0-:
-QAzphaQz71 RRRRRRRR-a-RERH#b8sFkRO0HDMOk#8CRV#F0sINCCR8PFCDbRC8L0$REzCRMCHPs0#H$VRF
A--zaQpQ1hz R7RRRRRR-R-RDBNHsVFM,HNRsAC	CCD$MRN80RH#FROMH0sLFk0s
#3-z-AQQpah z17RRRRRRRRR--ch3RCEH0C0sREMCRNRlCF0VREzCRMCHPs0#H$FRMsER0CNRMlRC#FHVR0-#
-QAzphaQz71 RRRRRRRR-O-RFsM0H0LkFRs#lRN$LkCR#RC80CFRMs8F#FCRssRbF0lFCsRbFO8k08#RCPsHC-8
-QAzphaQz71 RRRRRRRR-V-RsRFl0#EHRV#F0sINCHRI0kEF0bR#CVOHHbORssHFRHIs0M0CRsbCl#H#H3FM
A--zaQpQ1hz R7RRRRRR-R-
A--zaQpQ1hz R7RRRRRR-R-RQa]1mR1wqaW)Q R1)Rum7eQ A7RY]Ra  R)ta h1hRq7mRBhQa)Amza)`1R`Rq1Q'1'
A--zaQpQ1hz R7RRRRRR-R-R7qhRYqhRu X)1 1RRm)QpvuQR 7W)q)qQha R1,QphBzh7QtA,RzhaRmpaRQavQ a7Rm-,
-QAzphaQz71 RRRRRRRR-a-R]Q RvQup W7Rqq))h aQ1wRmR)v Bh]qaQqApYQaR7qhRawQh1 1R)wmR-q
-QAzphaQz71 RRRRRRRR-u-RqQ)aBqzp)zRu)1um )Rq QR71qBpQ7v 3hRQRRhm he a]R1qRppaR] )  thRa1m-)
-QAzphaQz71 RRRRRRRR-B-Rm)haQaAzmR)1Ap RQpqA mRw)hRqYQR7)a B,hRQ7 Q)BRa,QQhB7a hqRp,1Bu Q,qp
A--zaQpQ1hz R7RRRRRR-R-R  Xvqup)RY,mB)Rm h1Thz apQqRv7qq1t Rh5QB7pzQ,htRaAzRahmRvpQQ7a R,am
A--zaQpQ1hz R7RRRRRR-R-Rmu)B z)va hRRmw11zAazQaat Rm1m7RRm)1e )Q1B ;mRp1m1Rw1Rz 7,Rq,aqR
m)-z-AQQpah z17RRRRRRRRR--uw)mQ;a1RRm)AQz1h1 1RaQh z))umaQh]2RmeW  B)Rq z17hRq7hRmRYqhR a]m
)Y-z-AQQpah z17RRRRRRRRR--mpwRQQqApYQa,]RW  a])hRQRhBmaB)qa1,RaB)QaQRpqpAQQ,aYRRm)aam)
A--zaQpQ1hz R7RRRRRR-R-Rh5QB7pzQRhthp tQht Bm R)aRm]W )Q21 RQq)1tQhRRQhqRhYWRqYmRzamawR]- 
-QAzphaQz71 RRRRRRRR-z-R1m Rw]RaQ11RmWwaq,) R  ehwRQReq7Q71 RRmwaR] u1m1QpAQQRaYm1wRz
B]-z-AQQpah z17RRRRRRRRR--7qqvt
 3-z-AQQpah z17RRRRRRRR
---z-AQQpah z17RRRRRRRRR--h ma:ERaHe#R]R7pP#CsHRFMIRN#oCCMsCN08#RkHRMo0RECBCRPsF#HMVRFRC0E
A--zaQpQ1hz R7RRRRRR-R-RRRRRRRRRHFsoNHMDkRVMHO0FLMR$ER0C RQ e R]R7pvEN0C0lNHDONROuN	CNo
A--zaQpQ1hz R7RRRRRR-R-RRRRRRRRRsWF	oHMRFtsk5bRBK1/a-2
-QAzphaQz71 
A--zaQpQ1hz R7RRRRRRFROMN#0Mh0R:hRQa  t)=R:RU4.;-
-ApzQazQh1
 7-z-AQQpah z17RRRRRRRRR--aDNLCVRFRoDF52w[RD=RF_owE8CNrR[9+FRDo0w_NrHD[R9,VRFsw=[RR[4+/U4.3-
-ApzQazQh1R 7RRRRR-RR-#RzCV8RFosRCsMCNF0HMVRFR0CGCRM8bOsCHF#HMFRDoHNs0#El3-
-ApzQazQh1R 7RRRRR-RR-ERaCFROMN#0Md0R6c4Udj(.UdUU.#RHRc.^6#,RFER0CHR8PCH8RRH#COGN0-3
-QAzphaQz71 RRRRRRRR-Q-R0MRC#Cks#FROsOsC0CRsNM8HoVRFRoDFwC_ENR8,CMPCRsVFRNHMOsOkN
0C-z-AQQpah z17RRRRRRRRR--8HCOl-ND0LF-HsMN$FROMsPC#MHFRksF0CHM#53R sPC$8LF$CRo00#RE-C
-QAzphaQz71 RRRRRRRR-s-RH0oER#NMIRCsVRFsQ hat# )R#DC#ER0N.MR^36d2-
-ApzQazQh1R 7RRRRR-RR-NReD#kCRsVFRtpm5Rw2ICCsRMoCC0sNCk8R#oHMRsCsF<sRR^4j-R6(NFL#DCk0
A--zaQpQ1hz R7RRRRRR-R-R0IHEER0CORLRR-Db	NON3oC
A--zaQpQ1hz -7
-QAzphaQz71 RRRRRRRR0C$bRq) p _eB)amRRH#NNss$hR5q)azqspRNCMoR2<>RRFV)p q;-
-ApzQazQh1
 7-z-AQQpah z17RRRRRRRRMOF#M0N04Rq:q) p=R:Rjj3UddddddddddddU4(U;.(
A--zaQpQ1hz R7RRRRRRFROMN#0Mq0R. :)q:pR=3Rjj64.jjjjjdjj(((4cdg.;-
-ApzQazQh1R 7RRRRRORRF0M#NRM0q)d: Rqp:j=R3.jj.4d.dUgg(gg4cUc(j
g;-z-AQQpah z17RRRRRRRRMOF#M0N0cRq:q) p=R:Rjj3jdjcc(UU((((j4(ncc6(.-;
-QAzphaQz71 
A--zaQpQ1hz R7RRRRRRFROMN#0Mp0Rm_twapqQ: R)qep_ mBa)R5jahmR2=R:R-5
-QAzphaQz71 RRRRRRRRRRRRRRRRj,3j
A--zaQpQ1hz R7RRRRRRRRRRRRRRjR-3jjjjjjjjjjjj6jjc.d.gUgdcj.jc
g,-z-AQQpah z17RRRRRRRRRRRRRRRRjj3jjjjjjjjjjjjj.4((nc6(gcg(4jn,-
-ApzQazQh1R 7RRRRRRRRRRRRR-RRjj3jjjjjjjjjj4jjdj.d44(UUg...,dd
A--zaQpQ1hz R7RRRRRRRRRRRRRRjR-3jjjjjjjjjjjj4j46.c6(Un..UUg(
.,-z-AQQpah z17RRRRRRRRRRRRRRRR3-jjjjjjjjjjjjjjnjcng6.cgng6jUdj-,
-QAzphaQz71 RRRRRRRRRRRRRRRRjj3jjjjjjjjjj6jj4UcUc(g6.6nUU,4j
A--zaQpQ1hz R7RRRRRRRRRRRRRRjR-3jjjjjjjjjjjj6j.dn.4Udgc4c4(c
6,-z-AQQpah z17RRRRRRRRRRRRRRRR3-jjjjjjjjjjjjjj46.djn.n4dgdjn6c-,
-QAzphaQz71 RRRRRRRRRRRRRRRR-jj3jjjjjjjjjjjj4gU46jjnj4djn4UU,-
-ApzQazQh1R 7RRRRRRRRRRRRRjRR3jjjjjjjjjjjjdjn.ngj6Ug6(6.cc
c,-z-AQQpah z17RRRRRRRRRRRRRRRRjj3jjjjjjjjjjjjUcn46g4.dUnj(cU4,-
-ApzQazQh1R 7RRRRRRRRRRRRR-RRjj3jjjjjjjjjj(jjd(66(4j.g6cdj,.U
A--zaQpQ1hz R7RRRRRRRRRRRRRR3RjjjjjjjjjjjjjjdgnU(jnn66U6(..(-,
-QAzphaQz71 RRRRRRRRRRRRRRRRjj3jjjjjjjjjj(jj6ngUdgn6(c4g4,c4
A--zaQpQ1hz R7RRRRRRRRRRRRRR3Rjjjjjjjjjjjjjj(.6gggg4d.Ujgngj-,
-QAzphaQz71 RRRRRRRRRRRRRRRR-jj3jjjjjjjjjjjjccn6((.gcg(6Uccc,-
-ApzQazQh1R 7RRRRRRRRRRRRR-RRjj3jjjjjjjjjj(jj6g6n.Ujn(4c6d,dn
A--zaQpQ1hz R7RRRRRRRRRRRRRR3Rjjjjjjjjjjjjj4gj466(d.(.dj(Uc.-,
-QAzphaQz71 RRRRRRRRRRRRRRRR-jj3jjjjjjjjj4jj(gd4jcdcj.nc.ndj,-
-ApzQazQh1R 7RRRRRRRRRRRRR-RRjj3jjjjjjjjjj(jj(j4Ujd4dnUU.j,gU
A--zaQpQ1hz R7RRRRRRRRRRRRRR3Rjjjjjjjjjjjjj4Ujgjc(6jUgg6d6.U-,
-QAzphaQz71 RRRRRRRRRRRRRRRR-jj3jjjjjjjjjjjj.(jc.(d6Ucjjn64g,-
-ApzQazQh1R 7RRRRRRRRRRRRR-RRjj3jjjjjjjjjjUjjdj(.gg4jg6.dg,4.
A--zaQpQ1hz R7RRRRRRRRRRRRRR3Rjjjjjjjjjjjjj4UcjU(4.g4d(4d446-,
-QAzphaQz71 RRRRRRRRRRRRRRRRjj3jjjjjjjjjj.j4Ujng46(4(U6U.,6(
A--zaQpQ1hz R7RRRRRRRRRRRRRR3Rjjjjjjjjjjjjj4U((UjU6(4(UgjU4n-,
-QAzphaQz71 RRRRRRRRRRRRRRRRjj3jjjjjjjjjjnjjcUcj66n4jnngU,g4
A--zaQpQ1hz R7RRRRRRRRRRRRRR3Rjjjjjjjjjjjjj4dn4..U.n.n(c.jU.-,
-QAzphaQz71 RRRRRRRRRRRRRRRR-jj3jjjjjjjjjjjj(j6cg64n464gnU4U,-
-ApzQazQh1R 7RRRRRRRRRRRRR-RRjj3jjjjjjjjjjjjjj6dnjU(4U4Ud(,gj
A--zaQpQ1hz R7RRRRRRRRRRRRRR3Rjjjjjjjjjjjjjj.g4j(gd.gcg4Ucgc-,
-QAzphaQz71 RRRRRRRRRRRRRRRRjj3jjjjjjjjjjUj466n((6jggn(gj,4j
A--zaQpQ1hz R7RRRRRRRRRRRRRRjR-3jjjjjjjjjjjj4jdcng.66jn4cg4U
d,-z-AQQpah z17RRRRRRRRRRRRRRRR3-jjjjjjjjjjjjjjjgdggc6c4g6gUnUg-,
-QAzphaQz71 RRRRRRRRRRRRRRRRjj3jjjjjjjjjj(j4gd4cdjUn4gd.4,4(
A--zaQpQ1hz R7RRRRRRRRRRRRRRjR-3jjjjjjjjjjjjdj4j(.gg((4dUdjn
n,-z-AQQpah z17RRRRRRRRRRRRRRRRjj3jjjjjjjjj.jjd(jgd.U64U(6nggd,-
-ApzQazQh1R 7RRRRRRRRRRRRRjRR3jjjjjjjjjjjjg.dgcg6jccU.(44d
(,-z-AQQpah z17RRRRRRRRRRRRRRRRjj3jjjjjjjjj4jj6ddg(4(n(6cc6Ucj,-
-ApzQazQh1R 7RRRRRRRRRRRRR-RRjj3jjjjjjjjjjnjdUc(j.4Ud6(Udn,(U
A--zaQpQ1hz R7RRRRRRRRRRRRRR3Rjjjjjjjjjjjjjd.ngj6d(jjU.UUjjg-,
-QAzphaQz71 RRRRRRRRRRRRRRRR-jj3jjjjjjjjjjjjgddUc.4(.ndndgng,-
-ApzQazQh1R 7RRRRRRRRRRRRRjRR3jjjjjjjjjjjjcjgdgddUg4U6n4.g
j,-z-AQQpah z17RRRRRRRRRRRRRRRRjj3jjjjjjjjjcjj44cUd(4Uj6c.UU6n,-
-ApzQazQh1R 7RRRRRRRRRRRRR-RRjj3jjjjjjjjjjdjj(dg.4Uncjg.jd,4c
A--zaQpQ1hz R7RRRRRRRRRRRRRR3RjjjjjjjjjjjjjjjUcdn46d(jcg..cc-,
-QAzphaQz71 RRRRRRRRRRRRRRRR-jj3jjjjjjjjjdjjc..ngddccUU.6gc.,-
-ApzQazQh1R 7RRRRRRRRRRRRRjRR3jjjjjjjjjjjj(cd4g.44(g6c4.gc
6,-z-AQQpah z17RRRRRRRRRRRRRRRR3-jjjjjjjjjjjjj4(jc6j(6j(6U(cn64-,
-QAzphaQz71 RRRRRRRRRRRRRRRR-jj3jjjjjjjjj4jj4U44nd(4U6g6gdd.,-
-ApzQazQh1R 7RRRRRRRRRRRRRjRR3jjjjjjjjjjjj6d(c(g6((.6.U6g6
d,-z-AQQpah z17RRRRRRRRRRRRRRRRjj3jjjjjjjjj4jjd.g4U.c44g.4(66n,-
-ApzQazQh1R 7RRRRRRRRRRRRRjRR3jjjjjjjjjjjj(4j(c6(d(jd6n(.c
j,-z-AQQpah z17RRRRRRRRRRRRRRRRjj3jjjjjjjjj.jjg4dgU46gUc(nUjjj,-
-ApzQazQh1R 7RRRRRRRRRRRRR-RRjj3jjjjjjjjjj.jc(6gjjngjjjjn(,(c
A--zaQpQ1hz R7RRRRRRRRRRRRRR3Rjjjjjjjjjjjjj.(.(cnj(4j4cd6g66-,
-QAzphaQz71 RRRRRRRRRRRRRRRRjj3jjjjjjjjjjjj4U6cgn.gn.(gng,4.
A--zaQpQ1hz R7RRRRRRRRRRRRRRjR-3jjjjjjjjjjjjj.d(jdU46gc((j66
U,-z-AQQpah z17RRRRRRRRRRRRRRRRjj3jjjjjjjjj4jj64(n.(jd(ndgg6cd,-
-ApzQazQh1R 7RRRRRRRRRRRRRjRR3jjjjjjjjjjjjdjdc46(jg.n6jccU
.,-z-AQQpah z17RRRRRRRRRRRRRRRR3-jjjjjjjjjjjjjc.466U46jcndd.n4d-,
-QAzphaQz71 RRRRRRRRRRRRRRRRjj3jjjjjjjjjj.jdnn66ggUUn(gj4,cn
A--zaQpQ1hz R7RRRRRRRRRRRRRRjR-3jjjjjjjjjjjj(ccjnc.6jj4cc6.c
n,-z-AQQpah z17RRRRRRRRRRRRRRRRjj3jjjjjjjjjdjjc(6.ngc(6d.jg.((,-
-ApzQazQh1R 7RRRRRRRRRRRRR-RRjj3jjjjjjjjjj(jjjgcUng.d.g4j(,cn
A--zaQpQ1hz R7RRRRRRRRRRRRRR3Rjjjjjjjjjjjjj4(4(nUg((d64n4g.c-,
-QAzphaQz71 RRRRRRRRRRRRRRRR-jj3jjjjjjjjj4jjjc((dcc4nj4ngU6(,-
-ApzQazQh1R 7RRRRRRRRRRRRRjRR3jjjjjjjjjjjjU.4ncdddd.g.g464
j,-z-AQQpah z17RRRRRRRRRRRRRRRRjj3jjjjjjjjj.jjc.4dncdggd4dd44d,-
-ApzQazQh1R 7RRRRRRRRRRRRRjRR3jjjjjjjjjjjjjdg6n(c.g.jU(djj
j,-z-AQQpah z17RRRRRRRRRRRRRRRR3-jjjjjjjjjjjjj.(n6jgn(.6jdn6j(4-,
-QAzphaQz71 RRRRRRRRRRRRRRRRjj3jjjjjjjjjj(jd44d6c44gg.6gj,.4
A--zaQpQ1hz R7RRRRRRRRRRRRRRjR-3jjjjjjjjjjjj44(n.ng4nddjcU.d
4,-z-AQQpah z17RRRRRRRRRRRRRRRR3-jjjjjjjjjjjjj.6UnU6.U4g6(46cdd-,
-QAzphaQz71 RRRRRRRRRRRRRRRR-jj3jjjjjjjjj.jjd.U46.c.ncdcngUj,-
-ApzQazQh1R 7RRRRRRRRRRRRRjRR3jjjjjjjjjjjj6jn(6nngU(n6jUjn
.,-z-AQQpah z17RRRRRRRRRRRRRRRR3-jjjjjjjjjjjjj.4U.jd4cU4cnUn4.(-,
-QAzphaQz71 RRRRRRRRRRRRRRRRjj3jjjjjjjjjjjj4(gj4dn4(.c44.,6c
A--zaQpQ1hz R7RRRRRRRRRRRRRR3Rjjjjjjjjjjjjj44U4gndcdcnnc444j-,
-QAzphaQz71 RRRRRRRRRRRRRRRRjj3jjjjjjjjjjgjjUccjn(6.U..dn,.(
A--zaQpQ1hz R7RRRRRRRRRRRRRRjR-3jjjjjjjjjjjj4ddc6g4j..U(66.c
.,-z-AQQpah z17RRRRRRRRRRRRRRRR3-jjjjjjjjjjjjj4jUd.(U6dj6ncn4nU-,
-QAzphaQz71 RRRRRRRRRRRRRRRR-jj3jjjjjjjjj4jjn(.jc4jj6cn(cggc,-
-ApzQazQh1R 7RRRRRRRRRRRRRjRR3jjjjjjjjjjjjdcUj4ddcggc6.6dj
4,-z-AQQpah z17RRRRRRRRRRRRRRRR3-jjjjjjjjjjjjj(n46jd664d(.U4.46-,
-QAzphaQz71 RRRRRRRRRRRRRRRRjj3jjjjjjjjjjUjUU..4d4g6U46(U,66
A--zaQpQ1hz R7RRRRRRRRRRRRRRjR-3jjjjjjjjjjjjgdjjUj6jd64..dUc
c,-z-AQQpah z17RRRRRRRRRRRRRRRR3-jjjjjjjjjjjjjn(4jn466gU(.6g4cn-,
-QAzphaQz71 RRRRRRRRRRRRRRRRjj3jjjjjjjjjj6jdng6gnngnd(dcU,dj
A--zaQpQ1hz R7RRRRRRRRRRRRRR3RjjjjjjjjjjjjjdU6(.ndg6.g4(Undd-,
-QAzphaQz71 RRRRRRRRRRRRRRRR-jj3jjjjjjjjjcjjnn..jjU(jc46cU6(,-
-ApzQazQh1R 7RRRRRRRRRRRRRjRR3jjjjjjjjjjjj.n.(ng(.(g4.4.66
n,-z-AQQpah z17RRRRRRRRRRRRRRRRjj3jjjjjjjjj(jj.UUdg.c((n.j64(c,-
-ApzQazQh1R 7RRRRRRRRRRRRRjRR3jjjjjjjjjjjjU.njcgnn6n4.n44(
d,-z-AQQpah z17RRRRRRRRRRRRRRRR3-jjjjjjjjjjjjj4njgj6U.jjcn6(g.U-,
-QAzphaQz71 RRRRRRRRRRRRRRRRjj3jjjjjjjjjj.jjdg44cUgddjUj6,d(
A--zaQpQ1hz R7RRRRRRRRRRRRRRjR-3jjjjjjjjjjjjc6Un6gjU6jj..ggc
(,-z-AQQpah z17RRRRRRRRRRRRRRRR3-jjjjjjjjjjjjjjj.4dU(c.464cgccc-,
-QAzphaQz71 RRRRRRRRRRRRRRRR-jj3jjjjjjjjj.jjddd.4gU.cU66(Ucj,-
-ApzQazQh1R 7RRRRRRRRRRRRR-RRjj3jjjjjjjjjj.jcdnddgUc.U44cg,4n
A--zaQpQ1hz R7RRRRRRRRRRRRRRjR-3jjjjjjjjjjjjgcddddg(ggn(Ud(c
c,-z-AQQpah z17RRRRRRRRRRRRRRRRjj3jjjjjjjjjcjj44dcnjc((ddU666n,-
-ApzQazQh1R 7RRRRRRRRRRRRRjRR3jjjjjjjjjjjjUjncn4(d4nc6cg4n
n,-z-AQQpah z17RRRRRRRRRRRRRRRRjj3jjjjjjjjjcjj(66U6jdcjdccj4nc,-
-ApzQazQh1R 7RRRRRRRRRRRRRjRR3jjjjjjjjjjjjnUd((gnUcn((n6(g
6,-z-AQQpah z17RRRRRRRRRRRRRRRR3-jjjjjjjjjjjjjUn6(dc(dnncn6cUnj-,
-QAzphaQz71 RRRRRRRRRRRRRRRRjj3jjjjjjjjjj4j.g.4dU.4.gjdcj,g.
A--zaQpQ1hz R7RRRRRRRRRRRRRRjR-3jjjjjjjjjjjj.n.cc.U.n6dc4d4c
U,-z-AQQpah z17RRRRRRRRRRRRRRRR3-jjjjjjjjjjjjj4Ujgdc6gdc.6ddUcj-,
-QAzphaQz71 RRRRRRRRRRRRRRRRjj3jjjjjjjjjj6jndc4jd(4d(dndn,64
A--zaQpQ1hz R7RRRRRRRRRRRRRRjR-3jjjjjjjjjjjj6c(Ugj4g4j.((4jn
g,-z-AQQpah z17RRRRRRRRRRRRRRRR3-jjjjjjjjjjjjjd6(Uc4.6.cn66c(jj-,
-QAzphaQz71 RRRRRRRRRRRRRRRRjj3jjjjjjjjjjjjcg.dgd4d.UUn(n,nc
A--zaQpQ1hz R7RRRRRRRRRRRRRR3RjjjjjjjjjjjjjU.(ccddUgU4c6gU.4-,
-QAzphaQz71 RRRRRRRRRRRRRRRRjj3jjjjjjjjjj6j..44UU6Ucn.UcU,U.
A--zaQpQ1hz R7RRRRRRRRRRRRRRjR-3jjjjjjjjjjjjnjdjdU44jdnc6..6
(,-z-AQQpah z17RRRRRRRRRRRRRRRR3-jjjjjjjjjjjjj64j6U666g..cUjjg.-,
-QAzphaQz71 RRRRRRRRRRRRRRRRjj3jjjjjjjjjjUj(ncggj.ddd6d6d,4(
A--zaQpQ1hz R7RRRRRRRRRRRRRRjR-3jjjjjjjjjjjjjn(.(jUn4gngjcgn
j,-z-AQQpah z17RRRRRRRRRRRRRRRRjj3jjjjjjjjj4jjnU4j6((66ddg.Uc6,-
-ApzQazQh1R 7RRRRRRRRRRRRRjRR3jjjjjjjjjjjj66U.U(4Uncd.664j
g,-z-AQQpah z17RRRRRRRRRRRRRRRR3-jjjjjjjjjjjjjdc6.n((6.gg(jgc(4-,
-QAzphaQz71 RRRRRRRRRRRRRRRR-jj3jjjjjjjjj4jjU.d(jcUcg.6ngUj6,-
-ApzQazQh1R 7RRRRRRRRRRRRRjRR3jjjjjjjjjjjjnUUjUnngdU4cggc4
n,-z-AQQpah z17RRRRRRRRRRRRRRRRjj3jjjjjjjjjnjjnncU.jnU(n4cUj(j,-
-ApzQazQh1R 7RRRRRRRRRRRRRjRR3jjjjjjjjjjjjUndd44n6j4(n6cn4
g,-z-AQQpah z17RRRRRRRRRRRRRRRRjj3jjjjjjjjj.jj6c4c.(dj.(Udn.j(,-
-ApzQazQh1R 7RRRRRRRRRRRRR-RRjj3jjjjjjjjjj(j4.cdgc.c66cn4U2dc;-
-ApzQazQh1
 7-z-AQQpah z17RRRRRRRRMOF#M0N0mRpt]w_ :q7Rq) p _eB)am5ajRm2RhRR:=5-
-ApzQazQh1R 7RRRRRRRRRRRRRjRR3
j,-z-AQQpah z17RRRRRRRRRRRRRRRRjj3jU((.j4ccjc.nUjd4n.c,-
-ApzQazQh1R 7RRRRRRRRRRRRRjRR36j464jcUdn66dgn6n.ng
c,-z-AQQpah z17RRRRRRRRRRRRRRRRjj3.nd4(gj6.6U4cj(nUncj,-
-ApzQazQh1R 7RRRRRRRRRRRRRjRR3jjd(n(46nUnn6(n.nddc
(,-z-AQQpah z17RRRRRRRRRRRRRRRRjj3d4UdUcUnd4j.cn4.cUcU,-
-ApzQazQh1R 7RRRRRRRRRRRRRjRR36jcU6jgddnj4..c(n4c(
j,-z-AQQpah z17RRRRRRRRRRRRRRRRjj36cd.cc646U4Udj(nc666,-
-ApzQazQh1R 7RRRRRRRRRRRRRjRR3jjnnn.c.44UnncUg((UU
n,-z-AQQpah z17RRRRRRRRRRRRRRRRjj3n6(gj4nng6jU.c6gccc6,-
-ApzQazQh1R 7RRRRRRRRRRRRRjRR36j(.c.d.d4.(c6..jd6d
g,-z-AQQpah z17RRRRRRRRRRRRRRRRjj3Uc.cdgnn.g4jUcUcnU4d,-
-ApzQazQh1R 7RRRRRRRRRRRRRjRR3gjUn44.6UUngj(nndgj.
.,-z-AQQpah z17RRRRRRRRRRRRRRRRjj3g.n(gnn.cc6U6dc(4Un4,-
-ApzQazQh1R 7RRRRRRRRRRRRRjRR3d4j((gngUdn4(6n6c(Un
j,-z-AQQpah z17RRRRRRRRRRRRRRRR4j344jUcndnd.cjn4cdcd.j,-
-ApzQazQh1R 7RRRRRRRRRRRRRjRR3(44(jUdd66nnjcdjUj4d
n,-z-AQQpah z17RRRRRRRRRRRRRRRR4j3.jc(dUc(6jj4dj.U6jj(,-
-ApzQazQh1R 7RRRRRRRRRRRRRjRR344d6d(n6U((U(n4d.46d
n,-z-AQQpah z17RRRRRRRRRRRRRRRR4j3djUc..d.U.6gg..dngj.,-
-ApzQazQh1R 7RRRRRRRRRRRRRjRR364c4jU.jcgUc66(j.((g
6,-z-AQQpah z17RRRRRRRRRRRRRRRR4j3644gn.jcj(.6dn.4(j6d,-
-ApzQazQh1R 7RRRRRRRRRRRRRjRR3U46njj6d(j4ngn6jc6n6
4,-z-AQQpah z17RRRRRRRRRRRRRRRR4j3nc6.g.6(Udg6gUjUdn(U,-
-ApzQazQh1R 7RRRRRRRRRRRRRjRR344(U.6j6.ngnU64djc4n
j,-z-AQQpah z17RRRRRRRRRRRRRRRR4j3(jUc((n6cn(.Ujgnn(gc,-
-ApzQazQh1R 7RRRRRRRRRRRRRjRR3c4Ugd..dgUcdcUd44jc6
n,-z-AQQpah z17RRRRRRRRRRRRRRRR4j3gg4dc.U6g6ggnc6jn(jc,-
-ApzQazQh1R 7RRRRRRRRRRRRRjRR3(4gU(.6c.ddgU(6646.d
6,-z-AQQpah z17RRRRRRRRRRRRRRRR.j3j4c.646cc(.UnjndjUnn,-
-ApzQazQh1R 7RRRRRRRRRRRRRjRR3j.46(ncnjg4(jd6j(j.c
4,-z-AQQpah z17RRRRRRRRRRRRRRRR.j34(nUdUgdd6jj.6d4jn.c,-
-ApzQazQh1R 7RRRRRRRRRRRRRjRR3d..46cd644dccj.jjUj6
n,-z-AQQpah z17RRRRRRRRRRRRRRRR.j3.(gdc44jjUnc(.(d..nc,-
-ApzQazQh1R 7RRRRRRRRRRRRRjRR36.d6jnn(44d.jUnjnjd(
.,-z-AQQpah z17RRRRRRRRRRRRRRRR.j3c44(gngdUgUnn.njcU(6,-
-ApzQazQh1R 7RRRRRRRRRRRRRjRR3(.cU4dnnjdgcc6g.6Un(
(,-z-AQQpah z17RRRRRRRRRRRRRRRR.j364dg6g.jg(Ujd(.cj6.U,-
-ApzQazQh1R 7RRRRRRRRRRRRRjRR3g.6g66(.dccnnnUj6(4n
(,-z-AQQpah z17RRRRRRRRRRRRRRRR.j3nn6gdU6ccggnUjcjd(6(,-
-ApzQazQh1R 7RRRRRRRRRRRRRjRR34.(g(dd4U6ccjj4c4nd4
c,-z-AQQpah z17RRRRRRRRRRRRRRRR.j3(n(UU4c6jjjdUj(4.6cd,-
-ApzQazQh1R 7RRRRRRRRRRRRRjRR3d.U(4nU(dd4jU(dc6d.4
g,-z-AQQpah z17RRRRRRRRRRRRRRRR.j3Udgnd..g6gU.ccUd.nUg,-
-ApzQazQh1R 7RRRRRRRRRRRRRjRR36.gc.nc4g.Ud4c.j4ndg
g,-z-AQQpah z17RRRRRRRRRRRRRRRRdj3jn4.4jdd64(Ugjg(c(4(,-
-ApzQazQh1R 7RRRRRRRRRRRRRjRR3(djjj.6dg6.c(U.U6dj4
.,-z-AQQpah z17RRRRRRRRRRRRRRRRdj346.(6j(4j.jcd4g6(g(.,-
-ApzQazQh1R 7RRRRRRRRRRRRRjRR3Ud4c(6dd444U(jgcUgdg
j,-z-AQQpah z17RRRRRRRRRRRRRRRRdj3.4c4gUcnnd6c4dn(d46g,-
-ApzQazQh1R 7RRRRRRRRRRRRRjRR3gd.(.6dU(nd.g6(46nU.
U,-z-AQQpah z17RRRRRRRRRRRRRRRRdj3d66d646cg(.jnd.dcccU,-
-ApzQazQh1R 7RRRRRRRRRRRRRjRR3jdcg6.nU(ngjcc6jUU4g
.,-z-AQQpah z17RRRRRRRRRRRRRRRRdj3cnncn((nd4cnj.jUdUcU,-
-ApzQazQh1R 7RRRRRRRRRRRRRjRR34d6gc(n.6d4ncUU.jnnn
d,-z-AQQpah z17RRRRRRRRRRRRRRRRdj366(c6UUUg...d(4ngnd4,-
-ApzQazQh1R 7RRRRRRRRRRRRRjRR3.dngcj6gUdngj4c(d4.(
n,-z-AQQpah z17RRRRRRRRRRRRRRRRdj3n.Ud646n466Ug6g4(.d6,-
-ApzQazQh1R 7RRRRRRRRRRRRRjRR3dd((c4njgg(dcU4UU4Uc
j,-z-AQQpah z17RRRRRRRRRRRRRRRRdj3((gjU.d6gUdc4c4Undd6,-
-ApzQazQh1R 7RRRRRRRRRRRRRjRR3cdUcn44g4UgjU.g6nU.d
.,-z-AQQpah z17RRRRRRRRRRRRRRRRdj3U4g(n4(64ccjcnjcc4g6,-
-ApzQazQh1R 7RRRRRRRRRRRRRjRR3cdggUgdjcU.j.6cc4.44
(,-z-AQQpah z17RRRRRRRRRRRRRRRRcj3jcj.dc4n4c.(6cg(gg6(,-
-ApzQazQh1R 7RRRRRRRRRRRRRjRR36cjc4n6jjU4(gU44cj6g
U,-z-AQQpah z17RRRRRRRRRRRRRRRRcj346jngcg.gdU6d(UU6U66,-
-ApzQazQh1R 7RRRRRRRRRRRRRjRR36c4UU.(gc64dd6g4Ug6.
6,-z-AQQpah z17RRRRRRRRRRRRRRRRcj3.njggc.gn.ccd((dgd6c,-
-ApzQazQh1R 7RRRRRRRRRRRRRjRR3nc.jdUcg46dj4nUcn.gg
4,-z-AQQpah z17RRRRRRRRRRRRRRRRcj3d(44dccnU44Ud4jjcccn,-
-ApzQazQh1R 7RRRRRRRRRRRRRjRR3ncd.(dnn(n(c(6.c(g6.
n,-z-AQQpah z17RRRRRRRRRRRRRRRRcj3c(4.cj6nU4j6cdjgn4.U,-
-ApzQazQh1R 7RRRRRRRRRRRRRjRR3ncc.4U(j..nUUjc44nj4
d,-z-AQQpah z17RRRRRRRRRRRRRRRRcj36(4.ccnc4ndgd6j.cUd6,-
-ApzQazQh1R 7RRRRRRRRRRRRRjRR3nc6.cd(dUdc4cU(4.((d
.,-z-AQQpah z17RRRRRRRRRRRRRRRRcj3n(4466(44c..jgU.4j(g,-
-ApzQazQh1R 7RRRRRRRRRRRRRjRR3ncnj(Ug..ggcd6dcg6(n
j,-z-AQQpah z17RRRRRRRRRRRRRRRRcj3((jgg6(4.j4g(4d4d6gU,-
-ApzQazQh1R 7RRRRRRRRRRRRRjRR36c(Ugc6jncUgnU6Uggcc
(,-z-AQQpah z17RRRRRRRRRRRRRRRRcj3UUjnUg6.d6c6(4j(c..4,-
-ApzQazQh1R 7RRRRRRRRRRRRRjRR36cU6Uj(4U6(4.njc4jdc
g,-z-AQQpah z17RRRRRRRRRRRRRRRRcj3gjjddUgUj6c6..6dgdn6,-
-ApzQazQh1R 7RRRRRRRRRRRRRjRR36cgj.((ngn(Ucjd64cd(
4,-z-AQQpah z17RRRRRRRRRRRRRRRRcj3g.gU(gUn6n6n4j4cd.U.,-
-ApzQazQh1R 7RRRRRRRRRRRRRjRR3c6j6j6n46j(4.g4.g6dj
U,-z-AQQpah z17RRRRRRRRRRRRRRRR6j3jng.44gj(6gj.6d6.6dd,-
-ApzQazQh1R 7RRRRRRRRRRRRRjRR3d64g(c66j444ndc4cjcj
6,-z-AQQpah z17RRRRRRRRRRRRRRRR6j34jUn(c(n.djU6dcn(Ug6,-
-ApzQazQh1R 7RRRRRRRRRRRRRjRR3d6..4cUcnd(6U46njj.d
n,-z-AQQpah z17RRRRRRRRRRRRRRRR6j3.n(U(gjUnc.jUU6(6(c4,-
-ApzQazQh1R 7RRRRRRRRRRRRRjRR3.6dc(ncgnUUgc44jg4gj
U,-z-AQQpah z17RRRRRRRRRRRRRRRR6j3dc(j46cnUdg(c46g6ncd,-
-ApzQazQh1R 7RRRRRRRRRRRRRjRR346c6.g(Ud.c.44.6g(dc
(,-z-AQQpah z17RRRRRRRRRRRRRRRR6j3cdn4.(cd6cg(jn(.jggj,-
-ApzQazQh1R 7RRRRRRRRRRRRRjRR3j66n4c(46(g.cdg4(U.g
d,-z-AQQpah z17RRRRRRRRRRRRRRRR6j36c644(6j6ncj4j4.j6gn,-
-ApzQazQh1R 7RRRRRRRRRRRRRjRR3g66n(46Ud(g6gdg6(nn(
(,-z-AQQpah z17RRRRRRRRRRRRRRRR6j3n(cjjU4d.dU6U6(nn4n6,-
-ApzQazQh1R 7RRRRRRRRRRRRRjRR3U6n6(jcd66d.gnU(6cgn
4,-z-AQQpah z17RRRRRRRRRRRRRRRR6j3(4.ggd(66jn.4cU(j.g.,-
-ApzQazQh1R 7RRRRRRRRRRRRRjRR3(6(dd46nd6j6n.cg.c4n
j,-z-AQQpah z17RRRRRRRRRRRRRRRR6j3Ug4n4g(dnjd6n.4U4jgj,-
-ApzQazQh1R 7RRRRRRRRRRRRRjRR3n6Ujjcgcj6jdc4n(cg.d
d,-z-AQQpah z17RRRRRRRRRRRRRRRR6j3gUjd(nccn4j.j6(g(6jj,-
-ApzQazQh1R 7RRRRRRRRRRRRRjRR3c6g(4j(jc((nn.4g4dc(
c,-z-AQQpah z17RRRRRRRRRRRRRRRR6j3gjgjUg4Un.c6cjnn.c6g,-
-ApzQazQh1R 7RRRRRRRRRRRRRjRR3dnj.Ugj6d4cU4gcUnggU
(,-z-AQQpah z17RRRRRRRRRRRRRRRRnj3j6(66j.6.d.c.n.n.UnU,-
-ApzQazQh1R 7RRRRRRRRRRRRRjRR34n4U6j4cj44n6n4dgd46
6,-z-AQQpah z17RRRRRRRRRRRRRRRRnj34.njg(U(.n46.6dU6j6g,-
-ApzQazQh1R 7RRRRRRRRRRRRRjRR3jn..ccjj6g(4c.jc6.cd
(,-z-AQQpah z17RRRRRRRRRRRRRRRRnj3.dccdU.Ujd4.njgdd.jd,-
-ApzQazQh1R 7RRRRRRRRRRRRRjRR3Un.nnjU6.gc..(6n.Uj6
n,-z-AQQpah z17RRRRRRRRRRRRRRRRnj3dn.(ngnn6n(j.dUc(d.4,-
-ApzQazQh1R 7RRRRRRRRRRRRRjRR3nndgcj(nd..nc4gg(U(U
4,-z-AQQpah z17RRRRRRRRRRRRRRRRnj3cd4j4g4(cn.j(jg4g44(,-
-ApzQazQh1R 7RRRRRRRRRRRRRjRR36nc4gd(n(4ddjn.(gU.(
U,-z-AQQpah z17RRRRRRRRRRRRRRRRnj3c.g.(ngcnn.64j6jcjc6,-
-ApzQazQh1R 7RRRRRRRRRRRRRjRR3dn6d.j4(4.j4Ug6n(cc.
6,-z-AQQpah z17RRRRRRRRRRRRRRRRnj366(dU.j((jjgddj.U4g4,-
-ApzQazQh1R 7RRRRRRRRRRRRRjRR34nndcgUUc..6d.jg6..j
.,-z-AQQpah z17RRRRRRRRRRRRRRRRnj3n.6c..nd66ccj(64(6jn,-
-ApzQazQh1R 7RRRRRRRRRRRRRjRR3gnncndj6cdg.4gU(Udc(
4,-z-AQQpah z17RRRRRRRRRRRRRRRRnj3(.dc.6n(.d4.6cjc4.4c,-
-ApzQazQh1R 7RRRRRRRRRRRRRjRR3(n(dUgU.gd6jjg.jg(d4
4,-z-AQQpah z17RRRRRRRRRRRRRRRRnj3U64dgc..U.j(djU.n(.n,-
-ApzQazQh1R 7RRRRRRRRRRRRRjRR36nUdjjcjgdjU4.U4djjg
.,-z-AQQpah z17RRRRRRRRRRRRRRRRnj3Udg.d4.U.6dU6d(6U(j4,-
-ApzQazQh1R 7RRRRRRRRRRRRRjRR3dng44c(Unj6j(44(Ujdn;.2
A--zaQpQ1hz -7
-QAzphaQz71 RRRRRRRRPHNsNCLDRRv,Kh:Qa  t)-;
-QAzphaQz71 RRRRRRRRPHNsNCLDR,w4R,w.RRt,Tz,R,.Rz,:ReRq) p-;
-QAzphaQz71 RRRRRRRRPHNsNCLDR)Z m):R Rqp:j=R3-j;-8vNCNRPsLHND#CRFFRMRMOF#M0N0FRVDM8HoORFO#ks
A--zaQpQ1hz R7RRRRRRNRPsLHNDmCRhR :)p qRR:=4;3jRv--NR8CPHNsNCLDRR#FMOFRF0M#NRM0V8FDHRMoFkOOs-#
-QAzphaQz71 
A--zaQpQ1hz R7RRRRRR-R-Rk8FLRDCDLFo5R2,DG8Cb;52
A--zaQpQ1hz -7
-QAzphaQz71 RRRRRRRRPHNsNCLDR:z4)p q;-
-ApzQazQh1
 7-z-AQQpah z17RRRRCRLo
HM-z-AQQpah z17-
-ApzQazQh1R 7RRRRR-RR-ERBCRO	PHND8$H0RRFVNksol0CM
A--zaQpQ1hz R7RRRRRRVRHRX5RRR<=jR3j2ER0C-M
-QAzphaQz71 -$-#MC0E#RH#0MsN#0DNCV_FV-
-ApzQazQh1R 7RRRRRRRRRRRRRNRR#s#C0qRwp
1 -z-AQQpah z17RRRRRRRRRRRRRRRRRRRRRRRRbsCFRs0"<XR=3RjjMRHRtpm5"X2
A--zaQpQ1hz R7RRRRRRRRRRRRRRRRRRRRRRCR#PHCs0 $R)))m;-
-ApzQazQh1- 7-M#$0#ECH0#Rs#NMDCN0_
FM-z-AQQpah z17RRRRRRRRRRRRRRRR0sCk5sM)p q'Wpm2-;
-QAzphaQz71 RRRRRRRRCRM8H
V;-z-AQQpah z17-
-ApzQazQh1R 7RRRRR-RR-FRBl0bkCNRPDRkCVRFs#ObCHRNDOCN##-
-ApzQazQh1R 7RRRRRHRRVRR5XRR=4R3j2ER0C-M
-QAzphaQz71 RRRRRRRRRRRRRRRRskC0sjMR3
j;-z-AQQpah z17RRRRRRRR8CMR;HV
A--zaQpQ1hz -7
-QAzphaQz71 RRRRRRRRH5VRR=XRRavq]R_ 2ER0C-M
-QAzphaQz71 RRRRRRRRRRRRRRRRskC0s4MR3
j;-z-AQQpah z17RRRRRRRR8CMR;HV
A--zaQpQ1hz -7
-QAzphaQz71 RRRRRRRR-q-RslokCRM0skC8OF0HM4:RRR<=oRR<.G;R/l.^Ro=R;-
-ApzQazQh1R 7RRRRR-RR-RR$=*Rw5+4RRwV/2FRVsVR||=R<R-.^U-
-ApzQazQh1
 7-z-AQQpah z17RRRRRRRR:vR=pRQm5tAX
2;-z-AQQpah z17RRRRRRRR:tR=7Rp 5XuX-,Rv
2;-z-AQQpah z17RRRRRRRR:KR=hRQa  t) 5)qhp52t*5-j432R2;-B-RR8OFC8RN8j#R3V6RFssRF8kMH
Mo-z-AQQpah z17RRRRRRRRRw4:5=R4/3j)p q52h2R)*R 5qpK+2RRj43;-R-w44*.HUR#MRNRaQh )t RRHMrU4.,.649-
-ApzQazQh1R 7RRRRRwRR.=R:R-tRR;w4
A--zaQpQ1hz -7
-QAzphaQz71 RRRRRRRR-q-RbFbsGNHl0CCRGMbN#MHFRsVFRoDF5V4+.4/w2=R~R+kRR-J
-QAzphaQz71 RRRRRRRRt=R:Rj43/35.j4*w+2w.;-
-ApzQazQh1R 7RRRRRzRRRR:=.*3jwt.*;-
-ApzQazQh1R 7RRRRReRRRR:=z;*z
A--zaQpQ1hz R7RRRRRRRRT:z=R*5e*q+4RR5e*q+.RR5e*q+dRRqe*c222;-
-ApzQazQh1
 7-z-AQQpah z17RRRRRRRRR--BCN#RR4:k=4RRskRF8kMC08RF^R.-RcdNFL#DCk03HR1MROCkRR<.U^-,-
-ApzQazQh1R 7RRRRR-RR-RRRRRRRkE4RNN#R0FRl#d0R6HRL0R#,NRM8wk4*4#RHRNCGOR0,Nw#R4NRE#RR<UHRL0
#3-z-AQQpah z17RRRRRRRRR--RRRRR0RQR#NDF8RN8C#RG0NOD0$RFlR|*oDF.H_ERD+RFwo__NEC89r[R<|RRj(63-
-ApzQazQh1R 7RRRRR-RR--
-ApzQazQh1R 7RRRRRHRRVRR5K=R/RFjRsRRv/j=R2ER0C-M
-QAzphaQz71 RRRRRRRRRRRRRRRRz:4R=RRz+4R6d;3j
A--zaQpQ1hz R7RRRRRRRRRRRRRR4RzRR:=z-4RRd643
j;-z-AQQpah z17-
-ApzQazQh1R 7RRRRRRRRRRRRR-RR-NRB#.CR:4R|-RG|</R4.36nRCaERRl-NRM8[8-RCMbC80CMRs0ClN#RsxCRC
sF-z-AQQpah z17RRRRRRRRRRRRRRRRR--RRRRRkRR4RR=kFR0RR.cL#H03-
-ApzQazQh1R 7RRRRRRRRRRRRR-RR--
-ApzQazQh1R 7RRRRRCRRD
#C-z-AQQpah z17RRRRRRRRRRRRRRRRRz4:z=R;-
-ApzQazQh1R 7RRRRRRRRRRRRR-RR-za)hzB54R2;-M-QR0ORERH#Hk#R4RR=5k8FL2DCRD5VF2N0R45k2-
-ApzQazQh1R 7RRRRRCRRMH8RV-;
-QAzphaQz71 
A--zaQpQ1hz R7RRRRRR.RzRR:=5j.3*.5wRw-R44*z2RR-zw4*.*2RR
t;-z-AQQpah z17RRRRRRRRR--k+4RRRk.=VR./w5.+RV20CFRGN0sRCbsOHH#F
M3-z-AQQpah z17-
-ApzQazQh1R 7RRRRR-RR-FRDo25GRD=RF.o5^wl*44*5+/V.w242R-=
-QAzphaQz71 RRRRRRRR-5-RlF*DoE._Hm+pt]w_ 5q7[k2+4+2RR*5lD.Fo_+DFpwmt_Qaqp25[+;J2
A--zaQpQ1hz R7RRRRRR-R-RG5CN2O0R5+R0$HM2-
-ApzQazQh1
 7-z-AQQpah z17RRRRRRRRRz4:z=R4RR+)p q5*v2pwmt_q] 725hRp+Rm_tw]7 q5;K2RRRRRRRR- -RG0NO
A--zaQpQ1hz R7RRRRRR.RzRR:=5Rz.+mRptaw_q5QpKR22+;RTRRRRRRRR-a-RH
M$-z-AQQpah z17RRRRRRRRRz.:z=R.RR+pwmt_Qaqp25h*q) p25v;-
-ApzQazQh1R 7RRRRRsRRCs0kMzR54RR+z;.2
A--zaQpQ1hz R7RRMRC8mRpt
;

RRRRMVkOF0HMmRpt5.RXH:RM R)qRp2skC0s)MR RqpHR#
RRRRR-RR-CR7#HOsbF0HMR:
RRRRR-RR-RRRRRRRRC1CRMVkOF0HMCR8OsDNNF0HMMRHR Q  0R18jR4(.n3-g4gnR
RRRRRR-R-R0hFC
#:RRRRRRRR-R-RRRRRR2RNR0)Ck#sMRq) pm'pWMRFRsCsFRs
RLRRCMoH
RRRRRRRRR--BOEC	NRPDHH80F$RVsRNoCklM
0#RRRRRRRRH5VRR<XR=3RjjRR2RC0EM-
-#0$MEHC##sR0NDM#N_0CF
VVRRRRRRRRRRRRRRRRNC##sw0Rq p1
RRRRRRRRRRRRRRRRRRRRRRRRbsCFRs0"<XR=3RjjMRHRtpm.25X"R
RRRRRRRRRRRRRRRRRRRRRRCR#PHCs0 $R)))m;-
-#0$MEHC##sR0NDM#N_0CFRM
RRRRRRRRRRRRRsRRCs0kM 5)qpp'm;W2
RRRRRRRR8CMR;HV
R
RRRRRR-R-RlBFbCk0RDPNkVCRF#sRbHCONODRN##C
RRRRRRRRRHV5RRX=3R4jRR20MEC
RRRRRRRRRRRRRRRR0sCkRsMj;3j
RRRRRRRR8CMR;HV
R
RRRRRRVRHRX5RR.=R32jRRC0EMR
RRRRRRRRRRRRRRCRs0MksRj43;R
RRRRRRMRC8VRH;R

RRRRR-RR-FRBl0bkCNRPDRkCVRFsoCCMsRNDOCN#
RRRRRRRR0sCkRsM5qRvap]_m_t.m w_*tpm5RX22R;
RCRRMp8Rm;t.
R

RVRRk0MOHRFMp4mtjXR5:MRHRq) ps2RCs0kM R)qHpR#R
RRRRRR-R-R#7CObsH0MHF:R
RRRRRR-R-RRRRRRRR1RCCVOkM0MHFRO8CDNNs0MHFRRHMQ   R810R(4jn-3.4ngg
RRRRRRRRR--hCF0#R:
RRRRR-RR-RRRRRRRRRN2)kC0sRM#)p q'WpmRRFMCFsssR
RRCRLo
HMRRRRRRRR-B-RE	CORDPNH08H$VRFRoNskMlC0R#
RRRRRHRRVRR5X=R<Rjj3RR2R0MEC
#--$EM0C##HRN0sMN#D0FC_VRV
RRRRRRRRRRRRRRRRR#RN#0CsRpwq1R 
RRRRRRRRRRRRRRRRRRRRRsRRCsbF0XR"RR<=jR3jHpMRmjt45"X2
RRRRRRRRRRRRRRRRRRRRRRRRP#CC0sH$)R );m)
#--$EM0C##HRN0sMN#D0FC_MR
RRRRRRRRRRRRRRRRRR0sCk5sM)p q'Wpm2R;
RRRRRCRRMH8RV
;
RRRRRRRR-B-RFklb0PCRNCDkRsVFRC#bODHNR#ONCR#
RRRRRHRRVRR5XRR=4R3j2ER0CRM
RRRRRRRRRRRRRsRRCs0kM3RjjR;
RRRRRCRRMH8RV
;
RRRRRRRRH5VRR=XRR34jjRR20MEC
RRRRRRRRRRRRRRRR0sCkRsM4;3j
RRRRRRRR8CMR;HV
R
RRRRRR-R-RlBFbCk0RDPNkVCRFosRCsMCNODRN
#CRRRRRRRRskC0s5MRRavq]m_pt_4jm w_*tpm5RX22R;
RCRRMp8Rmjt4;


RRRRVOkM0MHFRtpmR:5XRRHM)p q;qRA1R :H)MR 2qpR0sCkRsM)p qR
H#RRRRRRRR-7-RCs#OHHb0F
M:RRRRRRRR-R-RRRRRRCR1CkRVMHO0F8MRCNODsHN0FHMRM RQ 1 R048Rj3(n.g-4gRn
RRRRR-RR-FRh0:C#
RRRRRRRRR--RRRRRNRR2CR)0Mks# R)qpp'mFWRMsRCs
FsRRRRLHCoMR
RRRRRR-R-RCBEOP	RN8DHHR0$FNVRslokC#M0
RRRRRRRRRHV5RRX<j=R32jRRER0C-M
-M#$0#ECH0#Rs#NMDCN0_VFV
RRRRRRRRRRRRRRRR#RN#0CsRpwq1R 
RRRRRRRRRRRRRRRRRRRRRsRRCsbF0XR"RR<=jR3jHpMRmXt5,qRA1" 2
RRRRRRRRRRRRRRRRRRRRRRRRP#CC0sH$)R );m)
#--$EM0C##HRN0sMN#D0FC_MR
RRRRRRRRRRRRRRsRRCs0kM 5)qpp'm;W2
RRRRRRRR8CMR;HV
R
RRRRRRVRHRA5RqR1 <j=R3FjRsqRA1= RRj43RR2R0MEC
RRRRRRRRRRRRRRRR#RN#0CsRpwq1R 
RRRRRRRRRRRRRRRRRRRRRsRRCsbF0AR"qR1 <j=R3FjRsqRA1= RRj43RRHMp5mtXA,Rq21 "R
RRRRRRRRRRRRRRRRRRRRRRCR#PHCs0 $R)))m;R
RRRRRRRRRRRRRRsRRCs0kM 5)qpp'm;W2
RRRRRRRR8CMR;HV
R
RRRRRR-R-RlBFbCk0RDPNkVCRF#sRbHCONODRN##C
RRRRRRRRRHV5RRX=3R4jRR20MEC
RRRRRRRRRRRRRRRR0sCkRsMj;3j
RRRRRRRR8CMR;HV
R
RRRRRRVRHRX5RRA=RqR1 2ER0CRM
RRRRRRRRRRRRRsRRCs0kM3R4jR;
RRRRRCRRMH8RV
;
RRRRRRRR-B-RFklb0PCRNCDkRsVFRMoCCDsNR#ONCR
RRRRRRCRs0MksRp5RmXt52m/ptq5A12 2;R
RRMRC8mRpt
;

R--RVRRk0MOHRFMRh1QRR5X:MRHRq) pRR2skC0s)MR RqpH-#
-RRRRRRRRR--7OC#s0HbH:FM
R--RRRRR-RR-RRRRRRRRCR1CkRVMHO0F8MRCNODsHN0FHMRM RQ 1 R048Rj3(n.g-4g-n
-RRRRRRRRR--hCF0#-:
-RRRRRRRRR--RRRRRRRRN12RQ-h5X=2RRQ-1h25X
R--RRRRR-RR-RRRRRRRR2RLRh1Q5RX2=RRXHqVRAX152RR< 
u1-R-RRRRRR-R-RRRRRRRRRRO215QhX=2RR-XRR*X*d!/dRRHV Ru1<ARq125XRA<Rq_1  
u1-R-RRRRRR-R-RRRRRRRRRR8215Qhv]qa__uQm)e _-.RRRX2=mRB125X
R--RRRRR-RR-RRRRRRRR2RCR1Bm5RX2=3R4jRR-j*36X.**RRHVq5A1X<2RR1 u
R--RRRRR-RR-RRRRRRRR2RVR1Bm5RX2=3R4jRR-j*36X.**R5+RXc**2!/cR
HV-R-RRRRRR-R-RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR1 u<ARq125XRq<A1  _u-1
--
-RRRRRRRRO#FM00NMR1 uR):R Rqp:A=Rq_1  *u1A q1_1 u;-R-RMBFPoCsCCMORHOs0HCsN-
-
R--RRRRRPRRNNsHLRDChRR:Q hat; )
R--RRRRRPRRNNsHLRDChq ta QeRA:Rm mpq:hR=RRX<3Rjj-;
-RRRRRRRRsPNHDNLCpRXmpBqR):R Rqp:q=RAX152
R;-R-RRRRRRNRPsLHNDeCRq pz: R)q
p;-R-RRRRRRNRPsLHNDaCR Rvu: R)q
p;---
-RRRRoLCH-M
-RRRRRRRRR--vCN	RmXpBRqp<qRva.]__
uQ-R-RRRRRRVRHRmXpBRqp>qRva.]__RuQ0MEC
R--RRRRRRRRRRRRRaRR Rvu:w=Rp)mm5mXpB/qpv]qa_u._Q
2;-R-RRRRRRRRRRRRRRpRXmpBqRR:=XBpmq-pRRva uq*va.]__;uQ
R--RRRRRCRRMH8RV-;
--
-RRRRRRRRHXVRpqmBpRR<jR3j0MEC
----M#$0#ECH0#Rs#NMDCN0_VFV
R--RRRRRRRRRRRRRNRR#s#C0qRwp
1 -R-RRRRRRRRRRRRRRRRRRRRRRCRsb0FsRp"XmpBqRR<=jR3jNCV0sCRs80kOHRFMH1MRQXh52-"
-RRRRRRRRRRRRRRRRRRRRRRRRP#CC0sH$)R );m)
----M#$0#ECH0#Rs#NMDCN0_
FM-R-RRRRRRRRRRRRRRpRXmpBqRR:=-mXpB;qp
R--RRRRRCRRMH8RV-;
--
-RRRRRRRR-B-RFklb0PCRNCDkRsVFRC#bODHNR#ONC-#
-RRRRRRRRRHVXBpmq=pRRjj3RsRFRmXpBRqp=qRva.]__RuQFXsRpqmBpRR=v]qa_RuQRC0EM-
-RRRRRRRRRRRRRRRRskC0sjMR3
j;-R-RRRRRRMRC8VRH;-
-
R--RRRRRHRRVXRRpqmBpRR=v]qa__uQm)e _0.RE
CM-R-RRRRRRRRRRRRRRVRHRth qeaQ ER0C-M
-RRRRRRRRRRRRRRRRRRRRRRRR0sCkRsM-j43;-
-RRRRRRRRRRRRRRRRCCD#
R--RRRRRRRRRRRRRRRRRRRRRsRRCs0kM3R4j-;
-RRRRRRRRRRRRRRRR8CMR;HV
R--RRRRRCRRMH8RV-;
--
-RRRRRRRRHRVRXBpmq=pRRavq]__dumQ_e_ ).ER0C-M
-RRRRRRRRRRRRRRRRRHVhq ta QeRC0EM-
-RRRRRRRRRRRRRRRRRRRRRRRRskC0s4MR3
j;-R-RRRRRRRRRRRRRRDRC#-C
-RRRRRRRRRRRRRRRRRRRRRRRR0sCkRsM-j43;-
-RRRRRRRRRRRRRRRRCRM8H
V;-R-RRRRRRMRC8VRH;-
-
R--RRRRRHRRVpRXmpBqR <Ru01RE
CM-R-RRRRRRRRRRRRRRVRHRth qeaQ ER0C-M
-RRRRRRRRRRRRRRRRRRRRRRRR0sCkRsM-mXpB;qp
R--RRRRRRRRRRRRRCRRD
#C-R-RRRRRRRRRRRRRRRRRRRRRRCRs0MksRmXpB;qp
R--RRRRRRRRRRRRRCRRMH8RV-;
-RRRRRRRR#CDC-
-RRRRRRRRRRRRRRRRHXVRpqmBpRR<A q1_1 uRC0EM-
-RRRRRRRRRRRRRRRRRRRRRRRRau vRR:=XBpmq-pRRp5XmpBq*mXpB*qpXBpmq/p2n;3j
R--RRRRRRRRRRRRRRRRRRRRRHRRV RhtQqae0 RE
CM-R-RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRCRs0MksR -av
u;-R-RRRRRRRRRRRRRRRRRRRRRRDRC#-C
-RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR0sCkRsMau v;-
-RRRRRRRRRRRRRRRRRRRRRRRRCRM8H
V;-R-RRRRRRRRRRRRRRMRC8VRH;-
-RRRRRRRRCRM8H
V;---
-RRRRRRRRva u=R:Ravq]Q_uRX-RpqmBp-;
-RRRRRRRRRHVq5A1au v2RR< Ru10MEC
R--RRRRRRRRRRRRRHRRV RhtQqae0 RE
CM-R-RRRRRRRRRRRRRRRRRRRRRRCRs0MksR -av
u;-R-RRRRRRRRRRRRRRDRC#-C
-RRRRRRRRRRRRRRRRRRRRRRRR0sCkRsMau v;-
-RRRRRRRRRRRRRRRRCRM8H
V;-R-RRRRRRDRC#-C
-RRRRRRRRRRRRRRRRRHVq5A1au v2RR<A q1_1 uRC0EM-
-RRRRRRRRRRRRRRRRRRRRRRRRau vRR:=au vR5-Rau v*va u *av/u2n;3j
R--RRRRRRRRRRRRRRRRRRRRRHRRV RhtQqae0 RE
CM-R-RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRCRs0MksR -av
u;-R-RRRRRRRRRRRRRRRRRRRRRRDRC#-C
-RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR0sCkRsMau v;-
-RRRRRRRRRRRRRRRRRRRRRRRRCRM8H
V;-R-RRRRRRRRRRRRRRMRC8VRH;-
-RRRRRRRRCRM8H
V;---
-RRRRRRRRva u=R:Ravq]__.u-QRRmXpB;qp
R--RRRRRHRRVARq1 5avRu2<uR 1ER0C-M
-RRRRRRRRRRRRRRRRRHVhq ta QeRC0EM-
-RRRRRRRRRRRRRRRRRRRRRRRRskC0saMR ;vu
R--RRRRRRRRRRRRRCRRD
#C-R-RRRRRRRRRRRRRRRRRRRRRRCRs0MksR -av
u;-R-RRRRRRRRRRRRRRMRC8VRH;-
-RRRRRRRRCCD#
R--RRRRRRRRRRRRRHRRVARq1 5avRu2<qRA1  _u01RE
CM-R-RRRRRRRRRRRRRRRRRRRRRR Rav:uR= Rav-uRR 5avau* *vuau v23/nj-;
-RRRRRRRRRRRRRRRRRRRRRRRRRHVhq ta QeRC0EM-
-RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRskC0saMR ;vu
R--RRRRRRRRRRRRRRRRRRRRRCRRD
#C-R-RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRCRs0MksR -av
u;-R-RRRRRRRRRRRRRRRRRRRRRRMRC8VRH;-
-RRRRRRRRRRRRRRRRCRM8H
V;-R-RRRRRRMRC8VRH;-
-
R--RRRRRaRR Rvu:q=RAv15q_a]umQ_e_ ).RR-XBpmq;p2
R--RRRRRHRRV Rav<uRR1 uRC0EM-
-RRRRRRRRRRRRRRRRau vRR:=4R3j- Ravau* *vuj;36
R--RRRRRRRRRRRRRHRRV RhtQqae0 RE
CM-R-RRRRRRRRRRRRRRRRRRRRRRCRs0MksR -av
u;-R-RRRRRRRRRRRRRRDRC#-C
-RRRRRRRRRRRRRRRRRRRRRRRR0sCkRsMau v;-
-RRRRRRRRRRRRRRRRCRM8H
V;-R-RRRRRRDRC#-C
-RRRRRRRRRRRRRRRRRHVau vRA<Rq_1  Ru10MEC
R--RRRRRRRRRRRRRRRRRRRRRaRR Rvu:4=R3-jRau v*va u3*j6RR+au v*va u *avau* /vu.jc3;-
-RRRRRRRRRRRRRRRRRRRRRRRRHhVR atqQRe 0MEC
R--RRRRRRRRRRRRRRRRRRRRRRRRRRRRRsRRCs0kMaR- ;vu
R--RRRRRRRRRRRRRRRRRRRRRCRRD
#C-R-RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRCRs0MksRva u-;
-RRRRRRRRRRRRRRRRRRRRRRRR8CMR;HV
R--RRRRRRRRRRRRRCRRMH8RV-;
-RRRRRRRR8CMR;HV

---R-RRRRRR Rav:uR=ARq1q5vad]___uQm)e _-.RRmXpB2qp;-
-RRRRRRRRHaVR Rvu<uR 1ER0C-M
-RRRRRRRRRRRRRRRRva u=R:Rj43Ra-R *vuau v*6j3;-
-RRRRRRRRRRRRRRRRHhVR atqQRe 0MEC
R--RRRRRRRRRRRRRRRRRRRRRsRRCs0kM Rav
u;-R-RRRRRRRRRRRRRRDRC#-C
-RRRRRRRRRRRRRRRRRRRRRRRR0sCkRsM-va u-;
-RRRRRRRRRRRRRRRR8CMR;HV
R--RRRRRCRRD
#C-R-RRRRRRRRRRRRRRVRHRva uRR<A q1_1 uRC0EM-
-RRRRRRRRRRRRRRRRRRRRRRRRau vRR:=4R3j-va u *avju*3+6RRva u *avau* *vuau v/3.cj-;
-RRRRRRRRRRRRRRRRRRRRRRRRRHVhq ta QeRC0EM-
-RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRskC0saMR ;vu
R--RRRRRRRRRRRRRRRRRRRRRCRRD
#C-R-RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRCRs0MksR -av
u;-R-RRRRRRRRRRRRRRRRRRRRRRMRC8VRH;-
-RRRRRRRRRRRRRRRRCRM8H
V;-R-RRRRRRMRC8VRH;-
-
R--RRRRR-RR-FRBl0bkCNRPDRkCVRFsoCCMsRNDOCN##-
-RRRRRRRRH5VR5mXpBRqp<qRvau]_Qe_m .)_RN2RM58RXBpmq>pRRjj3202RE
CM-S-SSeSRq pz:P=R_sOF8_HOlCF8_0sFNF0HMi5RBj,R3Rj,G.,R(4,R2-;
-RRRRRRRRRRRRRRRR-R-Rpeqz= :RmRB)B7Q5BRi,3RjjG,R,(R.,mR)aQqam5h24
2;-R-RRRRRRMRC8VRH;-
-
R--RRRRRhRRRR:=Q hatR )5pRwm5m)XBpmqvp/q_a]umQ_e_ ).;22
R--RRRRRORRNR#CT7zq)aqh5RRhlRF8cH2R#-
-RRRRRRRRRIRRERCMj>R=
S--SeSSq pz:P=R_sOF8_HOlCF8_0sFNF0HMi5RBj,R3Rj,XBpmqRp,.R(,4
2;-R-RRRRRRRRRRRRRR-R-ezqp =R:R)Bm75QBR,iBRjj3,pRXmpBq,(R.,mR)aQqam5h24
2;-R-RRRRRRRRRRCIEMRR4=->
-SSSSpeqz= :ROP_FHs8OF_l8sC_F00NH5FMR,iBRjj3,pRXmpBqRv-Rq_a]umQ_e_ )..,R(j,R2-;
-RRRRRRRRRRRRRRRRe--q pzRR:=B7m)QRB5iRB,j,3jRmXpBRqp-qRvau]_Qe_m .)_,(R.,-
-RRRRRRRRRRRRRRRR-R-RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRmR)aQqam5h2j
2;-R-RRRRRRRRRRCIEMRR.=->
-SSSSpeqz= :R_-PO8FsHlO_F_8CsNF00MHF5BRi,3RjjX,RpqmBpRR-v]qa_,uQR,.(R;42
R--RRRRRRRRRRRRR-RR-peqz: R=BR-mQ)7Bi5RBj,R3Rj,XBpmq-pRRavq]Q_u,(R.,mR)aQqam5h24
2;-R-RRRRRRRRRRCIEMRRd=->
-RSSRSRSezqp R:=-OP_FHs8OF_l8sC_F00NH5FMR,iBRjj3,pRXmpBqRv-Rq_a]dQ_u_ me),_.R,.(R;j2
R--RRRRRRRRRRRRR-RR-peqz: R=BR-mQ)7Bi5RBj,R3Rj,XBpmq-pRRavq]__dumQ_e_ )..,R(-,
-RRRRRRRRRRRRRRRRR--RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR)RRmaaqQ2mh5;j2
R--RRRRRCRRMO8RN;#C

---R-RRRRRRVRHRth qeaQ ER0C-M
-RRRRRRRRRRRRRRRR0sCkRsM-peqz
 ;-R-RRRRRRDRC#-C
-RRRRRRRRRRRRRRRR0sCkRsMezqp -;
-RRRRRRRR8CMR;HV
R--RCRRM18RQ
h;
-
-RVRRk0MOHRFMBRm15:XRRRHM)p q2CRs0MksRq) p#RH
R--RRRRR-RR-CR7#HOsbF0HM-:
-RRRRRRRRR--RRRRR1RRCVCRk0MOHRFM8DCON0sNHRFMHQMR R  1R084nj(34.-g
gn-R-RRRRRR-R-R0hFC
#:-R-RRRRRR-R-RRRRRRRRNB2Rm-15X=2RR1Bm5
X2-R-RRRRRR-R-RRRRRRRRLB2RmX152RR=15Qhv]qa__uQm)e _-.RR
X2-R-RRRRRR-R-RRRRRRRROB2Rmv15q_a]u+QRRRX2R-=RB5m1X-2
-RRRRRRRRR--RRRRR8RR2mRB125XR4=R3-jRRXX*/j.3RRHVq5A1X<2RR1 u
R--RRRRR-RR-RRRRRRRRRC2B5m1X=2RRj43Rj-R3X6**R*.+XR5*2*c/Rc!H-V
-RRRRRRRRR--RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRuR 1q<RAX152AR<q_1  
u1-R-RRRRRR-R-
R--RRRRRORRF0M#NRM0 Ru1: R)q:pR=qRA1  _uA1*q_1  ;u1

---R-RRRRRRNRPsLHNDXCRpqmBpRR:)p qRR:=q5A1X
2;-R-RRRRRRNRPsLHNDeCRq pz: R)q
p;-R-RRRRRRNRPsLHNDaCR Rvu: R)q
p;---
-RRRRoLCH-M
-RRRRRRRRR--vCN	RmXpBRqp<qRva.]__
uQ-R-RRRRRRVRHRmXpBRqp>qRva.]__RuQ0MEC
R--RRRRRRRRRRRRRaRR Rvu:w=Rp)mm5mXpB/qpv]qa_u._Q
2;-R-RRRRRRRRRRRRRRpRXmpBqRR:=XBpmq-pRRva uq*va.]__;uQ
R--RRRRRCRRMH8RV-;
--
-RRRRRRRRHXVRpqmBpRR<jR3j0MEC
----M#$0#ECH0#Rs#NMDCN0_VFV
R--RRRRRRRRRRRRRNRR#s#C0qRwp
1 -R-RRRRRRRRRRRRRRRRRRRRRRCRsb0FsRp"XmpBqRR<=jR3jNCV0sCRs80kOHRFMHBMRmX152-"
-RRRRRRRRRRRRRRRRRRRRRRRRP#CC0sH$)R );m)
----M#$0#ECH0#Rs#NMDCN0_
FM-R-RRRRRRRRRRRRRRpRXmpBqRR:=-mXpB;qp
R--RRRRRCRRMH8RV-;
--
-RRRRRRRR-B-RFklb0PCRNCDkRsVFRC#bODHNR#ONC-#
-RRRRRRRRRHVXBpmq=pRRjj3RsRFRmXpBRqp=qRva.]__RuQ0MEC
R--RRRRRRRRRRRRRsRRCs0kM3R4j-;
-RRRRRRRR8CMR;HV

---R-RRRRRRVRHRpRXmpBqRv=Rq_a]u0QRE
CM-R-RRRRRRRRRRRRRRCRs0MksR3-4j-;
-RRRRRRRR8CMR;HV

---R-RRRRRRVRHRmXpBRqp=qRvau]_Qe_m .)_RRFsXBpmq=pRRavq]__dumQ_e_ ).ER0C-M
-RRRRRRRRRRRRRRRR0sCkRsMj;3j
R--RRRRRCRRMH8RV-;
--
-RRRRRRRRau vRR:=q5A1XBpmq;p2
R--RRRRRHRRVRR5au vR <RuR120MEC
R--RRRRRRRRRRRRRsRRCs0kM4R53-jRR6j3*va u *av;u2
R--RRRRRCRRD
#C-R-RRRRRRRRRRRRRRVRHR 5av<uRR1Aq u_ 102RE
CM-R-RRRRRRRRRRRRRRRRRRRRRRCRs0MksR354jjR-3a6* *vuau vRa+R *vuau v*va u *av.u/c23j;-
-RRRRRRRRRRRRRRRRCRM8H
V;-R-RRRRRRMRC8VRH;-
-
R--RRRRRaRR Rvu:q=RAX15pqmBpvR-q_a].Q_u2-;
-RRRRRRRRRHV5 Rav<uRR1 u2ER0C-M
-RRRRRRRRRRRRRRRR0sCkRsM5j43Rj-R3a6* *vuau v2-;
-RRRRRRRR#CDC-
-RRRRRRRRRRRRRRRRH5VRau vRA<Rq_1  2u1RC0EM-
-RRRRRRRRRRRRRRRRRRRRRRRRskC0s5MR4R3j-6j3*va u *av+uRRva u *avau* *vuau v/3.cj
2;-R-RRRRRRRRRRRRRRMRC8VRH;-
-RRRRRRRRCRM8H
V;---
-RRRRRRRRva u=R:R1qARp5XmpBqRv-Rq_a]u;Q2
R--RRRRRHRRV Rav<uRR1 uRC0EM-
-RRRRRRRRRRRRRRRRskC0s5MR-j43Rj+R3a6* *vuau v2-;
-RRRRRRRR#CDC-
-RRRRRRRRRRRRRRRRH5VRau vRA<Rq_1  2u1RC0EM-
-RRRRRRRRRRRRRRRRRRRRRRRRskC0s5MR-j43R3+j6 *avau* Rvu- Ravau* *vuau v*va uc/.3;j2
R--RRRRRRRRRRRRRCRRMH8RV-;
-RRRRRRRR8CMR;HV

---R-RRRRRR-R-RlBFbCk0RDPNkVCRFosRCsMCNODRN##C
R--RRRRRsRRCs0kMQR1hq5vau]_Qe_m .)_RX-RpqmBp
2;-R-RR8CMR1Bm;R

RkRVMHO0FaMRq5hRXRR:H)MR 2qpR0sCkRsM)p qR
H#RRRRRRRR-7-RCs#OHHb0F
M:RRRRRRRR-R-RRRRRRCR1CkRVMHO0F8MRCNODsHN0FHMRM RQ 1 R048Rj3(n.g-4gRn
RRRRR-RR-FRh0:C#
RRRRRRRRR--RRRRRNRR2qRah35jj=2RRjj3
RRRRRRRRR--RRRRRLRR2qRahX5-2RR=-haq5
X2RRRRRRRR-R-RRRRRR2ROR0)Ck#sMRq) pm'pWMRFRsCsFHsRVRRX<3RjjR
RRRRRR-R-RRRRRRRR8)2RCs0kM)#R 'qp]]QtRRFMCFsssVRHR>XRRjj3
R
RRRRRRNRPsLHNDhCR atqQRe :mRAmqp h=R:R<XRRjj3;R
RRRRRRNRPsLHNDXCRpqmBpRR:)p qRR:=q5A1X;2R
RRRRRRRRsPNHDNLCqRep:z Rq) pR;
RRRRRPRRNNsHLRDCau vR):R ;qp
R
RRCRLo
HMRRRRRRRR-v-RNR	CjR3j<X=RpqmBp=R<Ravq]__.uRQ
RRRRRHRRVpRXmpBqRv>Rq_a].Q_uRC0EMR
RRRRRRRRRRRRRR Rav:uR=pRwm5m)XBpmqvp/q_a].Q_u2R;
RRRRRRRRRRRRRXRRpqmBp=R:RmXpBRqp- Ravvu*q_a].Q_u;R
RRRRRRMRC8VRH;R

RRRRRHRRVpRXmpBqRj<R30jRE
CM-$-#MC0E#RH#0MsN#0DNCV_FVR
RRRRRRRRRRRRRR#RN#0CsRpwq1R 
RRRRRRRRRRRRRRRRRRRRRsRRCsbF0XR"pqmBp=R<Rjj3R0NVCssRCO8k0MHFRRHMa5qhX
2"RRRRRRRRRRRRRRRRRRRRRRRR#CCPs$H0R) )m
);-$-#MC0E#RH#0MsN#0DNCM_F
RRRRRRRRRRRRRRRRmXpBRqp:-=RXBpmq
p;RRRRRRRRCRM8H
V;
RRRRRRRRR--BOEC	NRPDHH80F$RVsRNoCklMR0
RRRRRHRRVpRXmpBqRv=Rq_a]umQ_e_ ).ER0CRM
RRRRRRRRRRRRRNRR#s#C0qRwp
1 RRRRRRRRRRRRRRRRRRRRRRRRsFCbs"0RX#RHRlNRkHD0bRDCFvVRq_a]umQ_e_ ).MRHRhaq5"X2
RRRRRRRRRRRRRRRRRRRRRRRRP#CC0sH$)R );m)
RRRRRRRRRRRRRRRRRHVhq ta QeRC0EMR
RRRRRRRRRRRRRRRRRRRRRRCRs0Mks5q) pm'pW
2;RRRRRRRRRRRRRRRRCCD#
RRRRRRRRRRRRRRRRRRRRRRRR0sCk5sM)p q't]Q]
2;RRRRRRRRRRRRRRRRCRM8H
V;RRRRRRRRCRM8H
V;
RRRRRRRRRHVXBpmq=pRRavq]__dumQ_e_ ).ER0CRM
RRRRRRRRRRRRRNRR#s#C0qRwp
1 RRRRRRRRRRRRRRRRRRRRRRRRsFCbs"0RX#RHRlNRkHD0bRDCFvVRq_a]dQ_u_ me)R_.HaMRqXh52R"
RRRRRRRRRRRRRRRRRRRRR#RRCsPCHR0$ m)))R;
RRRRRRRRRRRRRHRRV RhtQqae0 RE
CMRRRRRRRRRRRRRRRRRRRRRRRRskC0s)M5 'qp]]Qt2R;
RRRRRRRRRRRRRCRRD
#CRRRRRRRRRRRRRRRRRRRRRRRRskC0s)M5 'qpp2mW;R
RRRRRRRRRRRRRRMRC8VRH;R
RRRRRRMRC8VRH;R

RRRRR-RR-FRBl0bkCNRPDRkCVRFs#ObCHRNDOCN##R
RRRRRRVRHRmXpBRqp=3RjjsRFRmXpBRqp=qRvau]_QER0CRM
RRRRRRRRRRRRRsRRCs0kM3RjjR;
RRRRRCRRMH8RV
;
RRRRRRRR-B-RFklb0PCRNCDkRsVFRMoCCDsNR#ONCR#
RRRRReRRq pzRR:=15QhXBpmq/p2B5m1XBpmq;p2
RRRRRRRRRHVhq ta QeRC0EMR
RRRRRRRRRRRRRRCRs0MksRq-ep;z 
RRRRRRRR#CDCR
RRRRRRRRRRRRRRCRs0MksRpeqz
 ;RRRRRRRRCRM8H
V;RCRRMa8Rq
h;
RRRVOkM0MHFRBq)1RQh5:XRRRHM)p qRs2RCs0kM R)qHpR#R
RRRRRR-R-R#7CObsH0MHF:R
RRRRRR-R-RRRRRRRR1RCCVOkM0MHFRO8CDNNs0MHFRRHMQ   R810R(4jn-3.4ngg
RRRRRRRRR--hCF0#R:
RRRRR-RR-RRRRRRRRRN2q1)BQ-h5X=2RR)-qBh1Q5
X2RRRRRRRR-R-RRRRRR2RLR0)Ck#sMRFXRMsRCs
Fs
RRRRRRRRsPNHDNLC RhtQqae: RRmAmph qRR:=XRR<j;3j
RRRRRRRRsPNHDNLCpRXmpBqR):R Rqp:q=RAX152R;
RRRRRPRRNNsHLRDCezqp RR:)p q;R

RCRLo
HMRRRRR-R-RCBEOP	RN8DHHR0$FNVRslokC#M0
RRRRHRRVpRXmpBqR4>R30jRE
CMRRRRRRRRR#N#CRs0w1qp R
RRRRRRRRRRRRRRCRsb0FsRA"q125XR4>R3HjRM)RqBh1Q5"X2
RRRRRRRRRRRRRRRRP#CC0sH$)R );m)
RRRRRRRRCRs0MksR
X;RRRRRMRC8VRH;R

RRRRRR--BbFlkR0CPkNDCFRVsbR#CNOHDNRO#
C#RRRRRVRHRmXpBRqp=3RjjER0CRM
RRRRRRRRskC0sjMR3
j;RRRRRDRC#RHVXBpmq=pRRj43RC0EMR
RRRRRRHRRV RhtQqae0 RE
CMRRRRRRRRRRRRRRRRskC0s-MRv]qa__uQm)e _
.;RRRRRRRRR#CDCR
RRRRRRRRRRRRRRCRs0MksRavq]Q_u_ me);_.
RRRRRRRRMRC8VRH;R
RRRRRCRM8H
V;
RRRR-RR-FRBl0bkCNRPDRkCVRFsoCCMsRNDOCN##R
RRRRRHXVRpqmBpRR<jR3g0MEC
RRRRRRRRqRepRz :q=R)qBahp5XmpBq/T51)4a53-jRRmXpB*qpXBpmq2p22R;
RRRRR#CDCR
RRRRRReRRq pzRR:=v]qa__uQm)e _-.RRBq)a5qh1aT)5j43RX-RpqmBpp*XmpBq2p/XmpBq2R;
RRRRR8CMR;HV
R
RRRRRHhVR atqQRe 0MEC
RRRRRRRRqRepRz :-=Rezqp R;
RRRRR8CMR;HV
R
RRRRRskC0seMRq pz;R
RR8CMRBq)1;Qh
R
RRMVkOF0HM)RqB1BmRR5X:MRHRq) ps2RCs0kM R)qHpR#R
RRRRRR-R-R#7CObsH0MHF:R
RRRRRR-R-RRRRRRRR1RCCVOkM0MHFRO8CDNNs0MHFRRHMQ   R810R(4jn-3.4ngg
RRRRRRRRR--hCF0#R:
RRRRR-RR-RRRRRRRRRN2qB)Bm-15X=2RRavq]Q_uRq-R)mBB125X
RRRRRRRRR--RRRRRLRR2CR)0Mks#RRXFCMRsssF
R
RRRRRRNRPsLHNDhCR atqQRe :mRAmqp h=R:R<XRRjj3;R
RRRRRRNRPsLHNDXCRpqmBpRR:)p qRR:=q5A1X
2;RRRRRRRRPHNsNCLDRpeqz: RRq) p
;
RLRRCMoH
RRRR-RR-ERBCRO	PHND8$H0RRFVNksol0CM
RRRRHRRVpRXmpBqR4>R30jRE
CMRRRRRRRRR#N#CRs0w1qp R
RRRRRRRRRRRRRRCRsb0FsRA"q125XR4>R3HjRM)RqB1Bm5"X2
RRRRRRRRRRRRRRRRP#CC0sH$)R );m)
RRRRRRRRCRs0MksR
X;RRRRRMRC8VRH;R

RRRRRR--BbFlkR0CPkNDCFRVsbR#CNOHDNRO#
C#RRRRRVRHR=XRRj43RC0EMR
RRRRRRsRRCs0kM3RjjR;
RRRRR#CDHXVRRj=R30jRE
CMRRRRRRRRR0sCkRsMv]qa__uQm)e _
.;RRRRRDRC#RHVXRR=-j43RC0EMR
RRRRRRsRRCs0kMqRvau]_QR;
RRRRR8CMR;HV
R
RRRRR-B-RFklb0PCRNCDkRsVFRMoCCDsNR#ONCR#
RRRRRRHVXBpmq>pRRgj3RC0EMR
RRRRRReRRq pzRR:=qa)Bq1h5T5)a4R3j-pRXmpBq*mXpB2qp/mXpB2qp;R
RRRRRCCD#
RRRRRRRRqRepRz :v=Rq_a]umQ_e_ ).RR-qa)BqXh5pqmBpT/1)4a53-jRRmXpB*qpXBpmq2p2;R
RRRRRCRM8H
V;
R
RRRRRHhVR atqQRe 0MEC
RRRRRRRRqRepRz :v=Rq_a]u-QRRpeqz
 ;RRRRRMRC8VRH;R

RRRRR0sCkRsMezqp R;
RMRC8)RqB1Bm;


RVRRk0MOHRFMqa)Bq5hRYRR:H)MR 2qpR0sCkRsM)p qR
H#RRRRRRRR-7-RCs#OHHb0F
M:RRRRRRRR-R-RRRRRRCR1CkRVMHO0F8MRCNODsHN0FHMRM RQ 1 R048Rj3(n.g-4gRn
RRRRR-RR-FRh0:C#
RRRRRRRRR--RRRRRNRR2)RqBhaq52-YR-=Rqa)BqYh52R
RRRRRR-R-RRRRRRRRLq2R)qBah25YR-=Rqa)Bq4h53Yj/2RR+v]qa__uQm)e _V.RF|sRY>|RRj43
RRRRRRRRR--RRRRRORR2)RqBhaq5RY2=RRYVRFs|RY|<uR 1R

RRRRRORRF0M#NRM0 Ru1: R)q:pR=qRA1  _uA1*q_1  *u1A q1_1 u;R

RRRRRPRRNNsHLRDChq ta QeRA:Rm mpq:hR=RRY<3RjjR;
RRRRRPRRNNsHLRDC)Q BuB)mq:pRRmAmph q;R
RRRRRRNRPsLHNDYCRpqmBpRR:)p qRR:=q5A1Y
2;RRRRRRRRPHNsNCLDRpeqz: RRq) p
;
RLRRCMoH
RRRR-RR-NRv	NCRslokCRM0|RY|<3=4jR
RRRRRHYVRpqmBpRR>4R3j0MEC
RRRRRRRRRRRRRRRRmYpBRqp:4=R3Yj/pqmBpR;
RRRRRRRRRRRRR)RR uBQ)qmBp=R:Rza) R;
RRRRR#CDCR
RRRRRRRRRRRRRR R)B)QumpBqRR:=w1qp R;
RRRRR8CMR;HV
R
RRRRR-B-RFklb0PCRNCDkRsVFRC#bODHNR#ONCR#
RRRRRRHVYBpmq=pRRjj3RC0EMR
RRRRRRHRRV R)B)QumpBqRC0EMR
RRRRRRRRRRRRRRVRHRth qeaQ ER0CRM
RRRRRRRRRRRRRRRRRRRRRsRRCs0kM-R5v]qa__uQm)e _;.2
RRRRRRRRRRRRRRRR#CDCR
RRRRRRRRRRRRRRRRRRRRRRCRs0MksRq5vau]_Qe_m .)_2R;
RRRRRRRRRRRRRCRRMH8RVR;
RRRRRRRRCCD#
RRRRRRRRRRRRRRRR0sCkRsMj;3j
RRRRRRRRMRC8VRH;R
RRRRRCRM8H
V;
RRRRHRRVpRYmpBqR <Ru01RE
CMRRRRRRRRRRHVhq ta QeRC0EMR
RRRRRRRRRRRRRRVRHRB) Qmu)BRqp0MEC
RRRRRRRRRRRRRRRRRRRRRRRR0sCkRsM5q-vau]_Qe_m .)_RY+RpqmBp
2;RRRRRRRRRRRRRRRRCCD#
RRRRRRRRRRRRRRRRRRRRRRRR0sCkRsM-mYpB;qp
RRRRRRRRRRRRRRRR8CMR;HV
RRRRRRRRDRC#RC
RRRRRRRRRRRRRHRRV R)B)QumpBqRC0EMR
RRRRRRRRRRRRRRRRRRRRRRCRs0MksRq5vau]_Qe_m .)_RY-RpqmBp
2;RRRRRRRRRRRRRRRRCCD#
RRRRRRRRRRRRRRRRRRRRRRRR0sCkRsMYBpmq
p;RRRRRRRRRRRRRRRRCRM8H
V;RRRRRRRRR8CMR;HV
RRRRCRRMH8RV
;
RRRRR-R-RlBFbCk0RDPNkVCRFosRCsMCNODRN##C
RRRReRRq pzRR:=R)Bm75QBRj43,pRYmpBq,3Rjj.,R(e,R mBa)tQhR.252
;
RRRRRVRHRB) Qmu)BRqp0MEC
RRRRRRRRqRepRz :v=Rq_a]umQ_e_ ).RR-ezqp R;
RRRRR8CMR;HV
R
RRRRRHhVR atqQRe 0MEC
RRRRRRRRpeqz: R=eR-q pz;R
RRRRRCRM8H
V;
RRRRsRRCs0kMqRep;z 
RRRCRM8qa)Bq
h;
R
RRMVkOF0HM)RqBhaqRR5Y:MRHRq) pX;RRH:RM R)qRp2skC0s)MR RqpHR#
RRRRR-RR-CR7#HOsbF0HMR:
RRRRR-RR-RRRRRRRRC1CRMVkOF0HMCR8OsDNNF0HMMRHR Q  0R18jR4(.n3-g4gnR
RRRRRR-R-R0hFC
#:RRRRRRRR-R-RRRRRRNRR2CR)0Mks#3RjjMRFRsCsF
s
RRRRRRRRPHNsNCLDRmYpBRqp: R)q
p;RRRRRRRRPHNsNCLDRpeqz: RRq) pR;
RCRLo
HM
RRRR-R-RCBEOP	RN8DHHR0$FNVRslokC#M0
RRRRVRHRR5Y=3RjjMRN8RRX=3RjjRR20MEC
RRRRRRRRRRRNC##sw0Rq p1RbsCF
s0RRRRRRRRRRRRRRRR"Bq)a5qhj,3jRjj32#RHR8kMCs0ClCHM8R"
RRRRRRRRRRRRR#RRCsPCHR0$ m)))R;
RRRRRRRRRCRs0MksRjj3;R
RRCRRMH8RV
;
RRRRRR--BbFlkR0CPkNDCFRVsbR#CNOHDNRO#
C#RRRRRRHVYRR=jR3j0MEC
RRRRRRRRRHVXRR>jR3j0MEC
RRRRRRRRRRRskC0sjMR3
j;RRRRRRRRCCD#
RRRRRRRRRRRskC0svMRq_a]u
Q;RRRRRRRRCRM8H
V;RRRRR8CMR;HV
R
RRHRRVRRX=3RjjER0CRM
RRRRRHRRVRRY>3RjjER0CRM
RRRRRRRRRCRs0MksRavq]Q_u_ me);_.
RRRRRRRR#CDCR
RRRRRRRRRR0sCkRsM-avq]Q_u_ me);_.
RRRRRRRR8CMR;HV
RRRRMRC8VRH;


RRRRRR--BbFlkR0CPkNDCFRVsCRoMNCsDNRO#
C#RRRRRmYpBRqp:q=RAY15/;X2
R
RReRRq pzRR:=qa)BqYh5pqmBp
2;
RRRRVRHR<XRRjj3RC0EMR
RRRRRReRRq pzRR:=v]qa_RuQ-qRep;z 
RRRRMRC8VRH;R

RRRRHYVRRj<R30jRE
CMRRRRRRRRRpeqz: R=eR-q pz;R
RRCRRMH8RV
;
RRRRR0sCkRsMezqp R;
RMRC8)RqBhaq;


RRRRVOkM0MHFRh1Q]XR5RH:RM R)qRp2skC0s)MR RqpHR#
RRRRR-RR-CR7#HOsbF0HMR:
RRRRR-RR-RRRRRRRRC1CRMVkOF0HMCR8OsDNNF0HMMRHR Q  0R18jR4(.n3-g4gnR
RRRRRR-R-R0hFC
#:RRRRRRRR-R-RRRRRR2RNR0)Ck#sMRX5 u25XR -RX-u5X/22.
3jRRRRRRRR-R-RRRRRR2RLRh1Q]X5-2RR=1]Qh5
X2
RRRRRRRRsPNHDNLC RhtQqae: RRmAmph qRR:=XRR<j;3j
RRRRRRRRsPNHDNLCpRXmpBqR):R Rqp:q=RAX152R;
RRRRRPRRNNsHLRDCau vR):R ;qp
RRRRRRRRsPNHDNLCqRepRz : R)q
p;
RRRRoLCHRM
RRRRR-RR-FRBl0bkCNRPDRkCVRFs#ObCHRNDOCN##R
RRRRRRVRHRmXpBRqp=3RjjER0CRM
RRRRRRRRRRRRRsRRCs0kM3RjjR;
RRRRRCRRMH8RV
;
RRRRRRRR-B-RFklb0PCRNCDkRsVFRMoCCDsNR#ONCR#
RRRRRaRR Rvu: =RXXu5pqmBp
2;RRRRRRRRezqp =R:R 5av-uRRj43/va uj2*3
6;
RRRRRRRRVRHRth qeaQ ER0CRM
RRRRRRRRRRRRReRRq pzRR:=-peqz
 ;RRRRRRRRCRM8H
V;
RRRRRRRR0sCkRsMezqp R;
RCRRM18RQ;h]
R
RRkRVMHO0FRMRB]m1RR5X:MRHRq) ps2RCs0kM R)qHpR#R
RRRRRR-R-R#7CObsH0MHF:R
RRRRRR-R-RRRRRRRR1RCCVOkM0MHFRO8CDNNs0MHFRRHMQ   R810R(4jn-3.4ngg
RRRRRRRRR--hCF0#R:
RRRRR-RR-RRRRRRRRRN2)kC0sRM#5u X5RX2+XR uX5-2.2/3Rj
RRRRR-RR-RRRRRRRRRL2B]m152-XRB=Rm51]X
2
RRRRRRRRPHNsNCLDRmXpBRqp: R)q:pR=ARq125X;R
RRRRRRNRPsLHNDaCR Rvu: R)q
p;RRRRRRRRPHNsNCLDRpeqz: RRq) pR;
RLRRCMoH
RRRRRRRRR--BbFlkR0CPkNDCFRVsbR#CNOHDNRO#
C#RRRRRRRRHXVRpqmBpRR=jR3j0MEC
RRRRRRRRRRRRRRRR0sCkRsM4;3j
RRRRRRRR8CMR;HV
R

RRRRR-RR-FRBl0bkCNRPDRkCVRFsoCCMsRNDOCN##R
RRRRRR Rav:uR=XR up5XmpBq2R;
RRRRReRRq pzRR:=5va uRR+4/3jau v23*j6
;
RRRRRRRRskC0seMRq pz;R
RRMRC8mRB1
];
RRRRMVkOF0HMaRRqRh]5:XRRRHM)p q2CRs0MksRq) p#RH
RRRRRRRRR--7OC#s0HbH:FM
RRRRRRRRR--RRRRR1RRCVCRk0MOHRFM8DCON0sNHRFMHQMR R  1R084nj(34.-g
gnRRRRRRRR-h-RF#0C:R
RRRRRR-R-RRRRRRRRN)2RCs0kM5#R 5XuX-2RRu X52-X2 /5XXu52RR+ 5Xu-2X2
RRRRRRRRR--RRRRRLRR2qRah-]5X=2RRq-ahX]52R

RRRRRPRRNNsHLRDChq ta QeRA:Rm mpq:hR=RRX<3RjjR;
RRRRRPRRNNsHLRDCXBpmq:pRRq) p=R:R1qA5;X2
RRRRRRRRsPNHDNLC Rav:uRRq) pR;
RRRRRPRRNNsHLRDCezqp RR:)p q;R

RLRRCMoH
RRRRRRRRR--BbFlkR0CPkNDCFRVsbR#CNOHDNRO#
C#RRRRRRRRHXVRpqmBpRR=jR3j0MEC
RRRRRRRRRRRRRRRR0sCkRsMj;3j
RRRRRRRR8CMR;HV
R
RRRRRR-R-RlBFbCk0RDPNkVCRFosRCsMCNODRN##C
RRRRRRRRva u=R:Ru X5mXpB2qp;R
RRRRRRqRepRz :5=Rau vR4-R3aj/ 2vu/ 5av+uRRj43/va u
2;
RRRRRRRRRHVhq ta QeRC0EMR
RRRRRRRRRRCRs0MksRq-ep;z 
RRRRRRRR#CDCR
RRRRRRRRRRCRs0MksRpeqz
 ;RRRRRRRRCRM8H
V;RRRRCRM8a]qh;R

RVRRk0MOHRFMq1)BQRh]5:XRRRHM)p q2CRs0MksRq) p#RH
RRRRRRRRR--7OC#s0HbH:FM
RRRRRRRRR--RRRRR1RRCVCRk0MOHRFM8DCON0sNHRFMHQMR R  1R084nj(34.-g
gnRRRRRRRR-h-RF#0C:R
RRRRRR-R-RRRRRRRRN)2RCs0kMp#RmRt5XRR+1aT)5*RXXRR+423j2R

RLRRCMoH
RRRRRRRRR--BbFlkR0CPkNDCFRVsbR#CNOHDNRO#
C#RRRRRRRRHXVRRj=R30jRE
CMRRRRRRRRRRRRRRRRskC0sjMR3
j;RRRRRRRRCRM8H
V;
RRRRRRRRR--BbFlkR0CPkNDCFRVsCRoMNCsDNRO#
C#RRRRRRRRskC0s5MRRtpm5RRX+TR1)Ra5XR*X+3R4jR222R;
RCRRMq8R)QB1h
];
R

RkRVMHO0FqMR)mBB15]RXRR:H)MR 2qpR0sCkRsM)p qR
H#RRRRRRRR-7-RCs#OHHb0F
M:RRRRRRRR-R-RRRRRRCR1CkRVMHO0F8MRCNODsHN0FHMRM RQ 1 R048Rj3(n.g-4gRn
RRRRR-RR-FRh0:C#
RRRRRRRRR--RRRRRNRR2CR)0Mks#mRptX5RR1+RT5)aRXX*R4-R32j2;RRRX=R>Rj43
RRRRRRRRR--RRRRRLRR2CR)0Mks#RRXFCMRsssF
R
RRCRLo
HMRRRRRRRR-B-RE	CORDPNH08H$VRFRoNskMlC0R#
RRRRRHRRVRRX<3R4jER0CRM
RRRRRRRRRRRRRRRRNC##sw0Rq p1
RRRRRRRRRRRRRRRRRRRRRRRRbsCFRs0"<XRRj43RRHMqB)Bm51]X
2"RRRRRRRRRRRRRRRRRRRRRRRR#CCPs$H0R) )m
);RRRRRRRRRRRRRRRRR0sCkRsMXR;
RRRRRCRRMH8RV
;
RRRRRRRR-B-RFklb0PCRNCDkRsVFRC#bODHNR#ONCR#
RRRRRHRRVRRX=3R4jER0CRM
RRRRRRRRRRRRRsRRCs0kM3RjjR;
RRRRRCRRMH8RV
;
RRRRRRRR-B-RFklb0PCRNCDkRsVFRMoCCDsNR#ONCR#
RRRRRsRRCs0kMRR5p5mtR+XRR)1TaX5R*-XRRj432;22
RRRR8CMRBq)B]m1;R

RVRRk0MOHRFMqa)BqRh]5:XRRRHM)p q2CRs0MksRq) p#RH
RRRRRRRRR--7OC#s0HbH:FM
RRRRRRRRR--RRRRR1RRCVCRk0MOHRFM8DCON0sNHRFMHQMR R  1R084nj(34.-g
gnRRRRRRRR-h-RF#0C:R
RRRRRR-R-RRRRRRRRN)2RCs0kM5#Rp5mtR354jRR+X52/4R3j-2RX2.2/3;jRRX|RR<|RRj43
RRRRRRRRR--RRRRRLRR2CR)0Mks#RRXFCMRsssF
RRRRoLCHRM
RRRRR-RR-ERBCRO	PHND8$H0RRFVNksol0CM#R
RRRRRRVRHR1qA5RX2>4=R30jRE
CMRRRRRRRRRRRRRRRRNC##sw0Rq p1
RRRRRRRRRRRRRRRRRRRRRRRRbsCFRs0"1qA5RX2>4=R3HjRM)RqBhaq]25X"R
RRRRRRRRRRRRRRRRRRRRRRCR#PHCs0 $R)))m;R
RRRRRRRRRRRRRRCRs0MksR
X;RRRRRRRRCRM8H
V;
RRRRRRRRR--BbFlkR0CPkNDCFRVsbR#CNOHDNRO#
C#RRRRRRRRHXVRRj=R30jRE
CMRRRRRRRRRRRRRRRRskC0sjMR3
j;RRRRRRRRCRM8H
V;
RRRRRRRRR--BbFlkR0CPkNDCFRVsCRoMNCsDNRO#
C#RRRRRRRRskC0sRM5j*36p5mtR354j2+X/354j2-XR22R;R
RRMRC8)RqBhaq]
;
CRM8Ravq] _)q
p;
