library verilog;
use verilog.vl_types.all;
entity cfg_cntl is
    generic(
        MASTER_SERI     : integer := 8;
        MASTER_PARA     : integer := 12;
        ASYNC_PERI      : integer := 13;
        SLAVE_SERI      : integer := 15;
        SLAVE_PARA      : integer := 9;
        FPSC_PARA       : integer := 7;
        MASTER_BYTE     : integer := 6;
        FLASH_SPI03     : integer := 5;
        FLASH_SPIX      : integer := 4;
        MPC_BYTE        : integer := 10;
        MPC_HWORD       : integer := 11;
        MPC_WORD        : integer := 14;
        CHK_PRE         : integer := 0;
        CHK_ID          : integer := 1;
        CHK_HDR         : integer := 2;
        CHK_FPGA        : integer := 3;
        CHK_RAM         : integer := 6;
        CHK_FPSC        : integer := 5;
        CHK_POST        : integer := 7;
        RESET_FSM       : integer := 0;
        CLR_RAM_FSM     : integer := 12;
        CFG_IDLE_FSM    : integer := 8;
        CONFIG_FSM      : integer := 24;
        ERR_IDLE_FSM    : integer := 9;
        USER_FSM        : integer := 26;
        PWRUP_BIT       : integer := 18
    );
    port(
        CCLK            : in     vl_logic;
        HCLK            : in     vl_logic;
        USR_START_CLK   : in     vl_logic;
        USR_GSR         : in     vl_logic;
        FPSC_GSR        : in     vl_logic;
        SYS_GSR         : in     vl_logic;
        RST_BUS         : in     vl_logic;
        RSTRAM          : in     vl_logic;
        GSRNRAM         : in     vl_logic;
        TRIRAM          : in     vl_logic;
        GSRN_SYNC_RAM   : in     vl_logic;
        RST_GSRN_RAM    : in     vl_logic;
        GSRN_INV_RAM    : in     vl_logic;
        SCLK_RAM        : in     vl_logic;
        DONE_RAM        : in     vl_logic_vector(1 downto 0);
        STRT_RAM        : in     vl_logic_vector(4 downto 0);
        TRI_RAM         : in     vl_logic_vector(3 downto 0);
        BS_MODE         : in     vl_logic;
        DONEIN          : in     vl_logic;
        INITIN_N        : in     vl_logic;
        CHK_STATE       : in     vl_logic_vector(2 downto 0);
        MATCH           : in     vl_logic;
        BAD_ADDR        : in     vl_logic;
        ERR_FLAG        : in     vl_logic_vector(1 downto 0);
        PTEST_N         : in     vl_logic;
        CFG_PRGM_N      : in     vl_logic;
        CFG_RESET_N     : in     vl_logic;
        AHB_DONE        : in     vl_logic;
        PRGM_JTAG       : in     vl_logic;
        PRGM_MPI        : in     vl_logic;
        PRGM_FPSC       : in     vl_logic;
        PRGM_USER       : in     vl_logic;
        EN_COUNT6       : in     vl_logic;
        OSC_DIV128      : in     vl_logic;
        PWRUP           : in     vl_logic;
        LMODE           : in     vl_logic_vector(3 downto 0);
        SYS_RST_RAM     : in     vl_logic;
        SYS_RST_N       : in     vl_logic;
        HRESET_OUT      : out    vl_logic;
        PAD_INIT_N      : out    vl_logic;
        FSM_RES_N       : out    vl_logic;
        FSM_INIT_RAM    : out    vl_logic;
        FSM_ERR         : out    vl_logic;
        PRGM_JTAG_N     : out    vl_logic;
        BS_RST_JTAG_N   : out    vl_logic;
        RST_LOCK        : out    vl_logic;
        PAD_DONE        : out    vl_logic;
        INIT_N          : out    vl_logic;
        TRI_ION         : out    vl_logic;
        DONE            : out    vl_logic;
        GSR_N           : out    vl_logic;
        GSRN_SYNC       : out    vl_logic;
        EN_PDWN         : out    vl_logic;
        PRGM_SYS        : out    vl_logic_vector(2 downto 0);
        PWR_ON          : out    vl_logic;
        PWRUPRES        : out    vl_logic
    );
end cfg_cntl;
