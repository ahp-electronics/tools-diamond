library verilog;
use verilog.vl_types.all;
entity PCNTR_sbnx8v1s is
    port(
        A               : in     vl_logic;
        Z               : out    vl_logic
    );
end PCNTR_sbnx8v1s;
