library verilog;
use verilog.vl_types.all;
entity config_register_func is
    port(
        edee            : in     vl_logic;
        xee             : in     vl_logic;
        all_dwnld_done  : in     vl_logic;
        refresh_out     : in     vl_logic;
        prog_128        : in     vl_logic;
        ext_done        : in     vl_logic;
        idcode          : in     vl_logic_vector(31 downto 0);
        clear_finish    : in     vl_logic;
        por             : in     vl_logic;
        tlreset         : in     vl_logic;
        tdi             : in     vl_logic;
        shiftir         : in     vl_logic;
        capir           : in     vl_logic;
        upir            : in     vl_logic;
        tck             : in     vl_logic;
        shiftdr         : in     vl_logic;
        updr            : in     vl_logic;
        capdr           : in     vl_logic;
        selbyp_b        : in     vl_logic;
        selbsr          : in     vl_logic;
        asrout_0        : in     vl_logic;
        dsrout_0        : in     vl_logic;
        bsout_0         : in     vl_logic;
        selasr          : in     vl_logic;
        mnfgshift       : in     vl_logic;
        idcode_o        : in     vl_logic;
        ucode_o         : in     vl_logic;
        ucode_ee_o      : in     vl_logic;
        progucode_sram_o: in     vl_logic;
        cmd_ld_ucode    : in     vl_logic;
        progdone_sram_o : in     vl_logic;
        progsec_sram_o  : in     vl_logic;
        progee_status   : in     vl_logic;
        readee_status   : in     vl_logic;
        flash_status    : in     vl_logic;
        flash_fail      : in     vl_logic;
        seldsr          : in     vl_logic;
        progdis_o       : in     vl_logic;
        progctrl0_o     : in     vl_logic;
        vfyctrl0_o      : in     vl_logic;
        cmd_prgm_done_r : in     vl_logic;
        cmd_prgm_done_comp: in     vl_logic;
        cmd_prgm_sec    : in     vl_logic;
        cmd_ld_ctrl0    : in     vl_logic;
        not_edit        : in     vl_logic;
        crc_err         : in     vl_logic;
        id_fail_r       : in     vl_logic;
        program         : in     vl_logic;
        erase_sram_o    : in     vl_logic;
        eraseall_sram_o : in     vl_logic;
        mux_clk         : in     vl_logic;
        wakeup          : in     vl_logic;
        cmd_ctrl0_r     : in     vl_logic_vector(31 downto 0);
        cmd_ucode_r     : in     vl_logic_vector(31 downto 0);
        seler1          : in     vl_logic;
        seler2          : in     vl_logic;
        er1out          : in     vl_logic;
        er2out          : in     vl_logic;
        jtag_unprogram  : in     vl_logic;
        jtag_functional : in     vl_logic;
        clear_memory    : in     vl_logic;
        selid           : in     vl_logic;
        edit_mod        : in     vl_logic;
        wakeup_clk      : in     vl_logic;
        rti             : in     vl_logic;
        cfg             : in     vl_logic_vector(1 downto 0);
        latch_shadow    : in     vl_logic;
        cfg_dd          : in     vl_logic;
        erase_pulse     : in     vl_logic;
        progsec_ee_o    : in     vl_logic;
        progdone_ee_o   : in     vl_logic;
        progcrc32_o     : in     vl_logic;
        read_crc_o      : in     vl_logic;
        read_crc_ee_o   : in     vl_logic;
        cmd_st_crc32    : in     vl_logic;
        chip_crc_2_reg  : in     vl_logic_vector(31 downto 0);
        ssi_en          : in     vl_logic;
        sso_en          : in     vl_logic;
        spisi           : in     vl_logic;
        sed_rdbk        : in     vl_logic;
        program_spi     : in     vl_logic;
        sspi_ucode_o    : in     vl_logic;
        sspi_ucode_ee_o : in     vl_logic;
        sspi_idcode_o   : in     vl_logic;
        sspi_vfyctrl0_o : in     vl_logic;
        sspi_vfyctrl0_ee_o: in     vl_logic;
        sspi_vfycrc32_o : in     vl_logic;
        sspi_vfycrc32_ee_o: in     vl_logic;
        sspi_progctrl0_ee_o: in     vl_logic;
        sspi_progucode_ee_o: in     vl_logic;
        sspi_progcrc32_ee_o: in     vl_logic;
        sspi_capdr      : in     vl_logic;
        progcrc32_ee_o  : in     vl_logic;
        progucode_ee_o  : in     vl_logic;
        nonjtag_cfg_r   : in     vl_logic;
        sed_enable_nedge: in     vl_logic;
        prem_time_out   : in     vl_logic;
        sospi           : in     vl_logic;
        status_out      : in     vl_logic;
        flash_mini      : in     vl_logic_vector(205 downto 0);
        flash_sec_l     : in     vl_logic_vector(3 downto 0);
        latch_encr      : in     vl_logic;
        sspi_refresh_o  : in     vl_logic;
        sspi_protect_o  : in     vl_logic;
        sspi_decrypt_o  : in     vl_logic;
        protect_shf_o   : in     vl_logic;
        decrypt_o       : in     vl_logic;
        dsrout_tag      : in     vl_logic;
        read_tag_o      : in     vl_logic;
        prog_tag_o      : in     vl_logic;
        sspi_read_tag_o : in     vl_logic;
        sspi_progsec_ee_o: in     vl_logic;
        sed_prgm_n      : in     vl_logic;
        cmd_crc         : in     vl_logic_vector(15 downto 0);
        read_crc16      : in     vl_logic;
        sspi_read_crc16 : in     vl_logic;
        sspi_rdstatus   : in     vl_logic;
        red_latch_rst   : in     vl_logic;
        sspi_progdis_o  : in     vl_logic;
        flclk           : in     vl_logic;
        refresh_o       : out    vl_logic;
        mclk_en_r       : out    vl_logic;
        mfgen           : out    vl_logic;
        mck_freq_switch : out    vl_logic;
        jtag_data       : out    vl_logic;
        jtag_addr       : out    vl_logic;
        instruction     : out    vl_logic_vector(7 downto 0);
        tdo_out         : out    vl_logic;
        tdo_en          : out    vl_logic;
        internal_done   : out    vl_logic;
        done_pupb       : out    vl_logic;
        freq_sel        : out    vl_logic_vector(5 downto 0);
        freq_div        : out    vl_logic_vector(5 downto 0);
        async_rst       : out    vl_logic;
        error           : out    vl_logic;
        done_reg        : out    vl_logic;
        program_effect  : out    vl_logic;
        init            : out    vl_logic;
        init_r          : out    vl_logic;
        mfg_bits        : out    vl_logic_vector(179 downto 0);
        e2_secty        : out    vl_logic;
        ues_crc_dsr     : out    vl_logic_vector(31 downto 0);
        done_ee_r       : out    vl_logic;
        auto_clear_en   : out    vl_logic;
        chip_crc_fm_reg : out    vl_logic_vector(31 downto 0);
        spi_prgm_clear  : out    vl_logic;
        sso             : out    vl_logic;
        freeze_io_en    : out    vl_logic;
        done_pin_override: out    vl_logic;
        done_pin_low    : out    vl_logic;
        status_cap      : out    vl_logic;
        status_shift    : out    vl_logic;
        encrypt_r       : out    vl_logic_vector(127 downto 0);
        key_r           : out    vl_logic;
        otp_active      : out    vl_logic;
        decrypt_en      : out    vl_logic;
        shf128_r        : out    vl_logic_vector(127 downto 0);
        sf_secty        : out    vl_logic;
        leave_postedit  : out    vl_logic
    );
end config_register_func;
