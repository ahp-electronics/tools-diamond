--
@ER--B$FbsEHo0OR52gR4g-cRRj.jd$R1MHbDO$H0ROQM
R--fN]C8:CsR#//$DMbH0OH$N/lb..jjDjdNl0/NCbbsN#/0D0/HoL/CFM_s6ONol/#k3D0PyE84
Rf-
-

R--****************************************************************R-R-
R--1MHoCv8RkHD0bCDHs-
-RsaNoRC0:NRp0O0HCsRmO6NR

---R-R4D3RFOoHRR-RNNss$kRlDb0HDsHCR0IHEHRbbkCLV5#RHOMRNR#CFbVRHDbCHMMHo-2
--R
-.RR3DRLFRO	-#RkHRMomNsORA6RD	FORDvk0DHbHRCs5pvzaX4U4
U2---
-BRRFsb$H0oER25ORj.jj.,RjRj41b$MDHHO0R$,Q3MO
R--RDqDRosHER0#sCC#s8PC3-
-
R--****************************************************************R-R-
-
-R****************************************************************-RR--
-RD#CCHO0F#MRC80RCMVHHF0HMR3R
R--NEsOD0H#RD=RFOoHRFLDOl	_k
D0-*-R*************************************************************R**R
--
R--****************************************************************R-R-
R--w#Hs0Fus80kO#,5qRRA,q
A2---
-HRW8q0ERI-RHE80RRFVqMRHb
k0-W-RHE80ARR-I0H8EVRFRHARM0bk
R--
R--q-ARR0LHI#NHChRq7VRFRDNDRbHMk
0#-
-R-*-R*************************************************************R**R
--
LDHs$NsRCHCC
;RkR#CHCCC38#0_oDFH4O_43ncN;DD
H
DLssN$sRFO;Nd
Ck#ROFsNFd3sOONF3lbN;DD
H
DLssN$$R#MHbDV
$;kR#C#b$MD$HV30N0skHL03C#N;DD
M
C0$H0RswH#s0uFO8k0H#R#R
RRMoCCOsH5R
RRRRRI0H8E:qRR0HMCsoC;R
RRRRRI0H8E:ARR0HMCsoC
RRR2R;
RFRbs50R
RRRRqRRRRR:HRMR#_08DHFoOC_POs0F58IH0-Eq4FR8IFM0R;j2
RRRRARRRRR:HRMR#_08DHFoOC_POs0F58IH0-EA4FR8IFM0R;j2
RRRRqRRARR:FRk0#_08DHFoOC_POs0F58IH0*EAI0H8E4q-RI8FMR0FjR2
RRRRRR--ARR*qR
RR
2;CRM8w#Hs0Fus80kO#
;
NEsOHO0C0CksRONsEF4RVHRwsu#0skF8OR0#H
#
R#RRHNoMD_RNNRkG:0R#8F_Do_HOP0COFIs5HE80qR-48MFI0jFR2R;
RHR#oDMNRNL_k:GRR8#0_oDFHPO_CFO0sH5I8A0E-84RF0IMF2Rj;C
Lo
HMRVRRFMsN8Rq:VRFsHHNRMRRj0IFRHE80qR-.oCCMsCN0
RRRRVRRFMsN8RA:VRFsHHLRMRRj0IFRHE80AR-.oCCMsCN0
RRRRRRRRARq58IH0*EAH+NRR2HLRR<=NN5H2MRN85RLH;L2
RRRRCRRMo8RCsMCNR0CVNFsM;8A
RRRRHRRVJ_C:VRHRN5HRj=R2CRoMNCs0RC
RRRRRRRRqIA5HE80A2-4RR<=N25jR8NMRIL5HE80A2-4;R
RRRRRCRM8oCCMsCN0R_HVC
J;RRRRRVRH_JMC:VRHRN5HRR/=jo2RCsMCN
0CRRRRRRRRR5qAI0H8EHA*NH+I8A0E-R42<5=RMRF0NN5H2N2RML8R58IH0-EA4
2;RRRRRMRC8CRoMNCs0HCRVC_MJR;
RMRC8CRoMNCs0VCRFMsN8
q;RVRRFMsN8RA:VRFsHHLRMRRj0IFRHE80AR-.oCCMsCN0
RRRRqRRAH5I8A0E*H5I8q0E-R42+LRH2=R<RIN5HE80q2-4R8NMRF5M05RLH2L2;R
RR8CMRMoCC0sNCFRVs8NMAR;
RRRRR5qAI0H8E5A*I0H8E4q-2RR+I0H8E4A-2=R<RIN5HE80q2-4R8NMRIL5HE80A2-4;M
C8sRNO;E4
-
-R****************************************************************-RR--
-R8N8s5CoqA,R,CR)#-2
--
-RPvFCs#RC#oH0#CsRR0FsDCbNROCbCHbL'kV#-
-R-
-R****************************************************************-RR-D

HNLssH$RC;CCR#
kCCRHC#C30D8_FOoH_n44cD3NDk;
#HCRC3CC#_08DHFoOM_k#MHoCN83D
D;
LDHs$NsROFsN
d;kR#CFNsOds3FOFNOlNb3D
D;
LDHs$NsRM#$bVDH$k;
##CR$DMbH3V$Ns00H0LkCN#3D
D;
0CMHR0$Ns88CHoR#R
RRMoCCOsH5R
RRRRRI0H8E:RRR0HMCsoC;R
RRRRRI0H8E:qRR0HMCsoC;R
RRRRRHCM8G:RRR0HMCsoC;R
RRRRRMLklC:sRR0HMCsoC;R
RRRRRsRCoR:RRR0HMCsoCRR--hCNlRRFV0RECDCCPDR
RR
2;RbRRFRs05R
RRRRRBRHM:MRHR8#0_oDFH
O;RRRRRRRqRRR:H#MR0D8_FOoH_OPC05FsI0H8ER-48MFI0jFR2R;
RRRRRRARRH:RM0R#8F_Do_HOP0COFIs5HE80-84RF0IMF2Rj;R
RRRRR)RC#:kRF00R#8F_Do_HOP0COFIs5HE80-84RF0IMF2Rj
RRR2R;
R0RN0LsHkR0C\N3sMR	\:MRH0CCosR;
R0RN0LsHkR0C\C3slCFP__MFIMNs\RR:HCM0o;Cs
8CMR8N8s;Co
s
NO0EHCkO0sNCRs4OERRFVNs88CHoR#R

RHR#oDMNR#)CkRD0:0R#8F_Do_HOP0COFIs5HE80-84RF0IMF2Rj;L

CMoH
RRR)kC#D<0R=RRq+RRA+HROMR;
RVRH_Rj:H5VRHCM8GRR>4o2RCsMCNR0C
RRRRVRRFFsDF:bjRsVFRHHRMRRj0IFRHE80qR-4oCCMsCN0
RRRRRRRR0RN0LsHkR0C\N3sMR	\FsVRCRo#:NRDLRCDHs#RC
o;RRRRRRRRR0N0skHL0\CR3lsCF_PCMIF_N\sMRRFVs#CoRD:RNDLCRRH#4R;
RRRRRoLCHRM
RRRRRRRRs#Co:HRbbkCLVR
RRRRRRRRRRFRbsl0RN
b5RRRRRRRRRRRRRRRRRRRQ=)>RCD#k025H,R
RRRRRRRRRRRRRRRRRm>R=R#)C5
H2RRRRRRRRRRRR2R;
RRRRR8CMRMoCC0sNCFRVsFDFb
j;RCRRMo8RCsMCNR0CR_HVj
;
RHRRV:_4RRHV58HMC=GRRR42oCCMsCN0RR
RRRRRVDFsF.Fb:FRVsRRHHjMRRR0FI0H8E4q-RMoCC0sNCR
RRRRRRNRR0H0sLCk0Rs\3N\M	RRFVs#CoqRR:DCNLD#RHRosC;R
RRRRRRNRR0H0sLCk0Rs\3CPlFCF_M_sINMF\RVCRsoR#q:NRDLRCDH4#R;R
RRRRRLHCoMR
RRRRRRsRRCqo#:HRbbkCLVR
RRRRRRRRRRFRbsl0RN
b5RRRRRRRRRRRRRRRRRRRQ=)>RCD#k025H,R
RRRRRRRRRRRRRRRRRm>R=R#)C5
H2RRRRRRRRRRRR2R;
RRRRR8CMRMoCC0sNCFRVsFDFb
.;RCRRMo8RCsMCNR0CR_HV4
;
RHRRV:_.RRHV5H.*MG8CRM=RkClLso2RCsMCNR0C
RRRRVRRFFsDF:bdRsVFRHHRMHRI8q0ERR0FI0H8ER-4oCCMsCN0
RRRRRRRR0RN0LsHkR0C\N3sMR	\FsVRCAo#RD:RNDLCRRH#s;Co
RRRRRRRR0RN0LsHkR0C\C3slCFP__MFIMNs\VRFRosC#:ARRLDNCHDR#;R4
RRRRLRRCMoH
RRRRRRRRCRso:#ARbbHCVLk
RRRRRRRRRRRRsbF0NRlbR5
RRRRRRRRRRRRRRRRR=QR>CR)#0kD5,H2
RRRRRRRRRRRRRRRRmRRRR=>)5C#HR2
RRRRRRRRR2RR;R
RRRRRCRM8oCCMsCN0RsVFDbFFdR;
RMRC8CRoMNCs0RCRH.V_;R

RVRH_Rd:H5VR.M*H8RCG<kRMlsLC2CRoMNCs0
CRRRRRRFRVsFDFbRc:VRFsHMRHR8IH0REq0IFRHE80-o4RCsMCN
0CRRRRRRRRR0N0skHL0\CR3MsN	F\RVCRsoR#B:NRDLRCDHs#RC
o;RRRRRRRRR0N0skHL0\CR3lsCF_PCMIF_N\sMRRFVs#CoBRR:DCNLD#RHR
4;RRRRRCRLo
HMRRRRRRRRRosC#RB:bCHbL
kVRRRRRRRRRRRRb0FsRblN5R
RRRRRRRRRRRRRRRRRQ>R=R#)Ck5D0H
2,RRRRRRRRRRRRRRRRRRRm=)>RCH#52R
RRRRRRRRRR;R2
RRRRCRRMo8RCsMCNR0CVDFsFcFb;R
RR8CMRMoCC0sNCHRRV;_d
8CMRONsE
4;
R--****************************************************************R-R-

---V-RDsFF5bQMkR0,mbk0k
02---
-*R**************************************************************R*R-
-
DsHLNRs$HCCC;kR
#HCRC3CC#_08DHFoO4_4nNc3D
D;kR#CHCCC38#0_oDFHNO_sEH03DND;#
kCCRHC#C30D8_FOoH_#kMHCoM8D3ND
;
DsHLNRs$FNsOdk;
#FCRsdON3OFsNlOFbD3ND
;
CHM00V$RDsFFR
H#RRRRRCRoMHCsO
R5RRRRRRRRRRRRI0H8ERQhRH:RMo0CC:sR=jRg;R
RRRRRRRRRRHRI8m0Ez:aRR0HMCsoCRR:=6
c;RRRRRRRRRRRRMLklCRsRRH:RMo0CC:sR=;R6
RRRRRRRRRRRR8IH0REqRRR:HCM0oRCs:6=R;R
RRRRRRRRRRMRH8RCGRRRR:MRH0CCos=R:4R
RRRRR2R;
RRRRRsbF0
R5RRRRRRRRRRRRQkMb0:RRRMRHR8#0_oDFHPO_CFO0sH5I8Q0EhR-48MFI0jFR2R;
RRRRRRRRRmRRkk0b0RR:FRk0#_08DHFoOC_POs0F58IH0zEmaR-48MFI0jFR2R
RRRRR2R;
RRRRR0N0skHL0\CR3MsN	:\RR0HMCsoC;R
SR0N0skHL0\CR3lsCF_PCMIF_N\sMRH:RMo0CC
s;CRM8VFDFs
;
NEsOHO0C0CksRONsEF4RVDRVFRFsH
#R
RRRRlOFbCFMMN0R8C8soR
RRoRRCsMCH5OR
RRRRRRRRHRI8R0ERH:RMo0CC
s;RRRRRRRRR8IH0REq:MRH0CCosR;
RRRRRRRRHCM8G:RRR0HMCsoC;R
RRRRRRMRRkClLsRR:HCM0o;Cs
RRRRRRRRCRsoRRRRH:RMo0CC-sR-NRhlFCRVER0CCRDP
CDRRRRR
2;RRRRRsbF0
R5RRRRRHRBMRR:H#MR0D8_FOoH;R
RRRRRqRRR:MRHR8#0_oDFHPO_CFO0sI5RHE80-84RF0IMF2Rj;R
RRRRRARRR:MRHR8#0_oDFHPO_CFO0sI5RHE80-84RF0IMF2Rj;R
RRRRR)RC#:kRF00R#8F_Do_HOP0COFIs5HE80-84RF0IMF2Rj
RRRR;R2
RRRCRM8ObFlFMMC0
;
R0RR$RbC#VEH0N_0LRDCHN#Rs$sNRk5MlsLC/8.RF0IMF2RjRRFVHCM0o;Cs
R
RRMVkOF0HMER#HxV0C5sFHCM8GRR:HCM0o2CsR0sCkRsM#VEH0N_0LRDCHR#
RRRRRsPNHDNLC0R#C:bRR0HMCsoC;R
RRRRRPHNsNCLDRL0NDPC_NRsR:ER#H_V00DNLCR;
RCRLo
HMRRRRR0R#C:bR=;R4
RRRRVRRFHsRRRHM4FR0R8HMC4G-RFDFbR
RRRRRR#RR0RCb:#=R0RCb*;R.
RRRRCRRMD8RF;Fb
RRRRVRRFHsRRRHMjFR0RlMkL/Cs.FRDFRb
RRRRRRRR0DNLCN_Ps25HRR:=#b0CR5*R.+*H4
2;RRRRRMRC8FRDF
b;RRRRRCRs0MksRL0NDPC_N
s;RCRRM#8RE0HVxFCs;R

RFROMN#0MD0RC0MoERR:HCM0oRCs:I=RHE80QMM/kClLsR;
RFROMN#0MI0RHE80ARR:HCM0oRCs:D=RC0MoERR-I0H8E
q;
RRRO#FM00NMRH#EV80N8RCs:ER#H_V00DNLC=R:RH#EVC0xsHF5MG8C2
;
LHCoMR
RRsVFDbFF_R4:VRFs[MRHR04RFkRMlsLC/o.RCsMCN
0CRLRRCMoH
RRRRsRRCqo#:8RN8osC
RRRRoRRCsMCHlORN5bR
RRRRIRRHE80RR=>DoCM0#E-E0HVNC88s-5[442-,R
RRRRRI0H8E=qR>HRI8q0E,R
RRRRRHCM8G>R=R
[,RRRRRkRMlsLCRR=>MLklC
s,RRRRRCRsoRRR=H>RMG8C
RRRR2RR
RRRRbRRFRs0l5Nb
RRRRRRRRRRRBRHM=Q>RM0bk5MDCo*0E5[.*-242,RR
RRRRRRRRq>R=RbQMkD05C0MoE.*5*4[-2R-48MFI0DFRC0MoE**.54[-2E+#HNV08s8C54[-22+4,R
RRRRRRARRRR=>QkMb0C5DMEo0*[.*-84RF0IMFCRDMEo0**5.[2-4+H#EV80N85Cs[2-4+,42
RRRRRRRRCR)#>R=R0mkb5k0DoCM0[E*-84RF0IMFCRDMEo0*-5[4#2+E0HVNC88s-5[442+2R
RRRRR2R;
RRRRRR--OsNs$FRVsER0CCRMGV0RDsFF
RRRRVRRFFsDFjb_:FRVsRRHHjMRRR0F#VEH08N8C[s5--42#VEH08N8Cjs52CRoMNCs0RC
RRRRRRRRRRRRRkRm00bk5MDCo*0E54[-2H+R2=R<R''j;R
RRRRRCRM8oCCMsCN0RsVFDbFF_
j;
RRRR-RR-DRNs8CN$CRoMNCs0
C8RRRRRFRVsFDFb:_NRsVFRHHRMRRj0#FRE0HVNC88s25j-o4RCsMCN
0CRRRRRRRRR0N0skHL0\CR3MsN	F\RVCRso:#RRLDNCHDR#MRH8;CG
RRRRRRRR0RN0LsHkR0C\C3slCFP__MFIMNs\VRFRosC#RR:DCNLD#RHR
4;RRRRRCRLo
HMRRRRRRRRRosC#b:RHLbCkRV
RRRRRRRRRRRRRFRbsl0RN
b5RRRRRRRRRRRRRRRRRRRRR=QR>MRQb5k0DoCM0.E**-5[4#2+E0HVNC88s-5[4#2-E0HVNC88s25j+H4+2R,
RRRRRRRRRRRRRRRRRRRRm>R=R0mkb5k0DoCM05E*[2-4+#H+E0HVNC88s-5[4#2-E0HVNC88s25j+
42RRRRRRRRRRRRRRRRRRRRR
2;RRRRRMRC8CRoMNCs0VCRFFsDFNb_;R

RMRC8CRoMNCs0VCRFFsDF4b_;R

RVRH_k#F#RN:H5VRMLklClsRF.8RR4=R2CRoMNCs0RC
RRRRR0N0skHL0\CR3MsN	F\RVCRsosONsR$#:NRDLRCDHH#RMG8C;R
RRRRRNs00H0LkC3R\sFClPMC_FN_IsRM\FsVRCNoOs#s$RD:RNDLCRRH#4R;
RCRLo
HMRRRRRFRVsFDFb:_dRsVFRHHRMRR40RFRDoCM0#E-E0HVNC88sk5MlsLC/-.24E+#HNV08s8C5Rj2oCCMsCN0
RRRRNRR0H0sLCk0Rs\3N\M	RRFVs#CoRD:RNDLCRRH#HCM8GR;
RRRRR0N0skHL0\CR3lsCF_PCMIF_N\sMRRFVs#CoRD:RNDLCRRH#4R;
RRRRRoLCHRM
RRRRRRRRs#Co:HRbbkCLVR
RRRRRRbRRFRs0l5Nb
RRRRRRRRRRRR=QR>MRQb5k0I0H8E-QhH
2,RRRRRRRRRRRRm>R=R0mkb5k0I0H8Eamz-
H2RRRRRRRRR
2;RRRRRMRC8CRoMNCs0VCRFFsDFdb_;R
RRRRRsOCoN$ss#b:RHLbCkRV
RRRRRRRRb0FsRblN5R
RRRRRRRRRRRRQ=Q>RM0bk58IH0hEQ-MDCo20E,R
RRRRRRRRRRRRm=m>Rkk0b0H5I8m0EzDa-C0MoER2
RRRRRRRR2R;
RRRRR0mkb5k0I0H8Eamz-MDCo+0E#VEH08N8CMs5kClLs2/.-H#EV80N85Csj82RF0IMFHRI8m0EzDa-C0MoE2+4RR<=
RRRRRRRRRRRRRRRQkMb0H5I8Q0EhC-DMEo0+H#EV80N85CsMLklC.s/2E-#HNV08s8C5Rj28MFI0IFRHE80QDh-C0MoE2+4;RR
RMRC8CRoMNCs0HCRVF_#k;#N
8CMRONsE
4;
LDHs$NsRCHCC
;RkR#CHCCC38#0_oDFH4O_43ncN;DD
Ck#RCHCC03#8F_Do_HON0sHED3NDk;
#HCRC3CC#_08DHFoOM_k#MHoCN83D
D;
LDHs$NsROFsN
d;kR#CFNsOds3FOFNOlNb3D
D;
0CMHR0$VFDFs8_N8RCsHR#
RRRRRMoCCOsHRR5
RRRRRRRRRIRRHE80QRhR:MRH0CCos=R:R;gj
RRRRRRRRRRRR8IH0zEmaRR:HCM0oRCs:6=RcR;
RRRRRRRRRMRRkClLsRRR:MRH0CCos=R:RR6
RRRRR
2;RRRRRFRbs50R
RRRRRRRRRRRRbQMkR0R:HRRM0R#8F_Do_HOP0COFIs5HE80Q4h-RI8FMR0Fj
2;RRRRRRRRRRRRmbk0k:0RR0FkR8#0_oDFHPO_CFO0sH5I8m0Ez4a-RI8FMR0FjR2
RRRRR
2;CRM8VFDFs8_N8;Cs
s
NO0EHCkO0sNCRs4OERRFVVFDFs8_N8RCsH
#RRORRF0M#NRM0DoCM0:ERR0HMCsoCRR:=I0H8E/QMMLklC
s;LHCoMR
RRsVFDbFF_R4:VRFs[MRHR04RFkRMlsLC/o.RCsMCN
0CRRRRRkRm00bk5MDCo*0E[R-48MFI0DFRC0MoE[*5-+424<2R=QRRM0bk5MDCo*0E5[.*--424FR8IFM0RMDCo*0E.[*5-+424R2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR+QkMb0C5DMEo0*[.*-84RF0IMFCRDMEo0**5.[2-4+
42RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR+RRRbQMkD05C0MoE.*5*4[-2
2;
RRRRmRRkk0b0C5DMEo0*-5[4R22<'=Rj
';RCRRMo8RCsMCNR0CVDFsF_Fb4
;
RHRRVF_#k:#NRRHV5lMkLRCslRF8.RR=4o2RCsMCN
0CRRRRRkRm00bk58IH0zEmaR-48MFI0IFRHE80m-zaDoCM0RE2<Q=RM0bk58IH0hEQ-84RF0IMFHRI8Q0EhC-DMEo02
;RRCRRMo8RCsMCNR0CH#V_FNk#;C

MN8Rs4OE;D

HNLssH$RC;CCR#
kCCRHC#C30D8_FOoH_n44cD3NDk;
#HCRC3CC#_08DHFoOs_NH30EN;DD
Ck#RCHCC03#8F_Do_HOkHM#o8MC3DND;C

M00H$8RN8aCss.CCR
H#RoRRCsMCH
O5RRRRRHRI8q0ERH:RMo0CC
s;RRRRRHRI8A0ERH:RMo0CC
s;RRRRRsR0CRCRRH:RMo0CCRs
R;R2
RRRb0FsRR5
RRRRRRq,qRl,ARR:H#MR0D8_FOoH;R
RRRRRqRAR:MRHR8#0_oDFHPO_CFO0sH5I8A0E*8IH0-Eq4FR8IFM0R;j2
RRRRbRRskF8O:0RR0FkR8#0_oDFHPO_CFO0sH5I8A0E+8IH0-Eq4FR8IFM0R
j2RRRRR-R-R*ARRRq
R;R2
8CMR8N8CssaC;C.
NR
sHOE00COkRsCNEsO4VRFR8N8CssaCRC.HR#
RFROMN#0M00REHCEo:ERR8#0_oDFHPO_CFO0s654RI8FMR0Fj:2R=mRBh1e_ap7_mBtQ_Be a5m)I0H8E4q-,nR42R;
RFROlMbFCRM0VFDFsR
RRRRRoCCMsRHO5R
RRRRRRIRRHE80QRhR:MRH0CCos
R;RRRRRRRRR8IH0zEmaRR:HCM0oRCs;R
RRRRRRMRRkClLsRRR:MRH0CCos
R;RRRRRRRRR8IH0REqRRR:HCM0oRCs;R
RRRRRRHRRMG8CRRRR:MRH0CCosR
RRRRR2R;
RRRRRFRbs50R
RRRRRRRRRRRRQRRM0bkRRR:H#MR0D8_FOoH_OPC05FsI0H8E-Qh4FR8IFM0R;j2
RRRRRRRRRRRRmRRkk0b0RR:FRk0#_08DHFoOC_POs0F58IH0zEmaR-48MFI0jFR2R
RRRRRR
2;RCRRMO8RFFlbM0CM;R

RFROlMbFCRM0VFDFs8_N8
CsRRRRRCRoMHCsO
R5RRRRRRRRR8IH0hEQRRR:HCM0oRCs;R
RRRRRRIRRHE80mRza:MRH0CCos
R;RRRRRRRRRlMkLRCsRRR:HCM0o
CsRRRRR;R2
RRRRRRRb0FsRR5
RRRRRRRRRRRRRbQMkR0R:MRHR8#0_oDFHPO_CFO0sH5I8Q0EhR-48MFI0jFR2R;
RRRRRRRRRRRRR0mkbRk0:kRF00R#8F_Do_HOP0COFIs5HE80m-za4FR8IFM0R
j2RRRRR2RR;R
RR8CMRlOFbCFMM
0;
RRRVOkM0MHFRb8C0HEW8R0EskC0sHMRMo0CCHsR#R
RRoLCHRM
RRRRVRFsHMRHRR468MFI0jFRRFDFbR
RRRHV5C0EEEHo5RH2=4R''02RE
CMRRRRRCRs0MksR4H+;R
RR8CMR;HV
RRRRMRC8FRDF
b;RRRRR0sCkRsMjR;
RMRC8CR8bW0EHE80;R

RFROMN#0M80RCEb0RH:RMo0CC:sR=CR8bW0EHE80;R
RRMOF#M0N0HRI800ERH:RMo0CC:sR=HRI8A0E+8IH0+Eq.R;
R$R0bDCRHRl#HN#Rs$sNRC58b+0E4FR8IFM0RRj2FHVRMo0CC
s;RR
RRMVkOF0HMNRODkOhlsLC#CRs0MksRlDH##RH
RRRRPRRNNsHLRDC0_ECMLklCRs#:HRDl
#;RLRRCMoH
RRRR0RREMC_kClLsj#52=R:R8IH0;Eq
RRRRVRRFHsRRRHM4FR0Rb8C04E+RFDFbR
RRRRRR0RREMC_kClLsH#52=R:RC0E_lMkL#Cs54H-2R/.+0R5EMC_kClLsH#5-R42lRF8.
2;RRRRRMRC8FRDF
b;RRRRRCRs0MksRC0E_lMkL#Cs;R
RRMRC8NRODkOhlsLC#R;

RRRO#FM00NMRlMkL#CsRD:RHRl#:O=RNhDOkClLs
#;RR
RRMVkOF0HMNRODHOplCRs0MksRlDH##RH
RRRRPRRNNsHLRDC0_ECD#HlRD:RH;l#
RRRRPRRNNsHLRDCMLklRH:RMo0CC
s;RLRRCMoH
RRRR0RREDC_H5l#j:2R=;Rj
RRRRMRRkRlL:I=RHE80qR;
RRRRRsVFRHHRMRR408FRCEb0+D4RF
FbR0RREDC_H5l#H:2R=ER0CH_DlH#5-R42+kRMlIL*HE800R;
RkRMl:LR=kRMl.L/R5+RMLklR8lFR;.2
RRRRCRRMD8RF;Fb
RRRRsRRCs0kMER0CH_Dl
#;RRRRCRM8OONDp;Hl
RR
RFROMN#0MP0RCHODlRR:D#HlRR:=OONDp;Hl
RRR#MHoNLDRHso0C:CRR8#0_oDFHPO_CFO0sC5POlDH5b8C04E+2R-48MFI0jFR2R;
RHR#oDMNRsONsR$,#MHo,HR#oRM4:0R#8F_Do;HO
C
LoRHM
RRRH	V_C_CbNC88sCasCH:RV0R5sRCC=2RjRMoCC0sNC-R-RCk#RsVFRbbHCMDHHRMoNRM8DRFIO0F#
R
RRRRR#MHoRR<=qFRGs;RA
RRRR#RRH4oMRR<=qsRFR
A;RRRRRNROsRs$<5=RMRF0qRl2NRM8AR;
RRRRRoLH0CsC58IH0-E04FR8IFM0RRj2<R=RBemh_71a_tpmQeB_ mBa),5jR8IH02Eq
RRRRRRRRRRRRRRRRRRRRRRRRRRRR&RRRsONsR$
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRq&RAH5I8A0E-84RF0IMF2Rj
RRRRRRRRRRRRRRRRRRRRRRRRRRRR&RRRhBmea_17m_pt_QBea Bmj)5,2R4;R

RRRRRsVFNqM8:FRVsNRHRRHM4FR0R8IH0-EqdCRoMNCs0RC
RRRRRRRRL0Hos5CC5+HN4I2*HE800R-48MFI0HFRNH*I800E2=R<RmRBh1e_ap7_mBtQ_Be a5m)jI,RHE80q-+4H
N2RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR&qIA5HE80AH*5N2+4-84RF0IMFHRI8A0E*2HN
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR&RRRhBmea_17m_pt_QBea Bmj)5,NRH+;42
RRRRCRRMo8RCsMCNR0CVNFsM;8q
RRRR-RR-MRFCCRLVCFsRC0ER#DN0CRPOs0F
RRRRLRRHso0C5C5I0H8E4q-2H*I800E-84RF0IMFIR5HE80q2-.*8IH02E0RR<=RhBmea_17m_pt_QBea Bmj)5,2R.
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR#&RH
oMRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR&ARq58IH0*EA58IH0-Eq442-RI8FMR0FI0H8E5A*I0H8E.q-2R2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR&RRRhBmea_17m_pt_QBea Bmj)5,HRI8q0E-;42
RRRR-RR-NRD#P0RCFO0sR
RRRRRL0Hos5CCI0H8EIq*HE800R-48MFI05FRI0H8E4q-2H*I800E2=R<RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRmRBh1e_ap7_mBtQ_Be a5m)j4,R2R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR&RRRo#HMR4
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR&ARq58IH0*EAI0H8E4q-RI8FMR0FI0H8E5A*I0H8E4q-2R2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR&mRBh1e_ap7_mBtQ_Be a5m)jI,RHE80q2-4
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR&q
;
RRRRRFRVsFDFbV.:F[sRRRHM4FR0Rb8C0oERCsMCN
0CRRRRRRRRR:l4RDRVF
FsRRRRRRRRRRRRoCCMsRHOlRNb5R
RRRRRRRRRRRRRRRRRRIRRHE80QRhR=P>RCHODl25[RP-RCHODl-5[4
2,RRRRRRRRRRRRRRRRRRRRR8IH0zEma>R=ROPCD5Hl[2+4RP-RCHODl25[,R
RRRRRRRRRRRRRRRRRRMRRkClLsRRR=M>RkClLs[#5-,42
RRRRRRRRRRRRRRRRRRRRHRI8q0ER=RR>HRI8q0E,R
RRRRRRRRRRRRRRRRRRHRRMG8CRRRR=[>R
RRRRRRRRRRRRR2
RRRRRRRRRbRRFRs0lRNb5R
RRRRRRRRRRRRRRRRRRQRRM0bkRRRR=L>RHso0CPC5CHODl25[-84RF0IMFCRPOlDH54[-2
2,RRRRRRRRRRRRRRRRRRRRR0mkbRk0R>R=RoLH0CsC5OPCD5Hl[2+4-84RF0IMFCRPOlDH52[2
RRRRRRRRRRRR
2;RRRRRMRC8oRRCsMCNR0CVDFsF.Fb;R
RR8CMRMoCC0sNCVRH_C	Cb8_N8aCss;CC
R
RR_HVM	F0C_CbNC88sCasCH:RV0R5sRCC=2R4RMoCC0sNC-R-RCk#RRHVNC88sVRN0RCs0RECl0kDHHbDCRs
RRRRRR--I0H8E>qR=
RcRRRRRHR#oRMR<q=RRsGFR
A;RRRRRHR#oRM4<q=RRRFsAR;
RRRRRsONs<$R=MR5Fq0RlN2RMA8R;R
RRRRRL0Hos5CCI0H8E40-RI8FMR0Fj<2R=BRRm_he1_a7pQmtB _eB)am5Rj,I0H8E
q2RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR&OsNs$R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRR&ARq58IH0-EA4FR8IFM0R
j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR&Bemh_71a_tpmQeB_ mBa),5jR;42
R
RRRRRHIV_HE80qH:RVIR5HE80qRR>do2RCsMCN
0CRRRRRRRRRoLH0CsC5I.*HE800R-48MFI0IFRHE800<2R=BRRm_he1_a7pQmtB _eB)am5Rj,I0H8E
q2RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR&RRR5qA.H*I8A0E-84RF0IMFHRI8A0E2R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRq&R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR&;Rq
R
RRRRRRVRRFMsN8Rq:VRFsHHNRMRR.0IFRHE80qR-doCCMsCN0
RRRRRRRRRRRRoLH0CsC5N5H+*42I0H8E40-RI8FMR0FHIN*HE800<2R=BRRm_he1_a7pQmtB _eB)am5Rj,I0H8E4q+-2HN
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR&qIA5HE80AH*5N2+4-84RF0IMFHRI8A0E*2HN
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR&qR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR&RRRhBmea_17m_pt_QBea Bmj)5,NRH2R;
RRRRRRRRCRM8oCCMsCN0RsVFNqM8;R
RRRRRR-RR-MRFCCRLVCFsRC0ER#DN0CRPOs0F
RRRRRRRRHRLoC0sCI55HE80q2-4*8IH0-E04FR8IFM0RH5I8q0E-*.2I0H8ER02<R=RBemh_71a_tpmQeB_ mBa),5jR
.2RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR&RRRo#HMR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRq&RAH5I8A0E*H5I8q0E--424FR8IFM0R8IH0*EA58IH0-Eq.
22RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR&RRRRq
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR&Bemh_71a_tpmQeB_ mBa),5jR8IH0-Eq.
2;RRRRRMRC8CRoMNCs0HCRVH_I8q0E;R

RRRRR_HVI0H8Ejq_:VRHRH5I8q0ERd=R2CRoMNCs0RC
RRRRRRRR-F-RMLCRCsVFCER0CNRD#P0RCFO0sR
RRRRRRLRRHso0C.C5*8IH0-E04FR8IFM0R8IH02E0RR<=RhBmea_17m_pt_QBea Bmj)5,2R.
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR&HR#oRM
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR&q.A5*8IH0-EA4FR8IFM0R8IH02EA
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR&
RqRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR&RRR
q;
RRRRCRRMo8RCsMCNR0CHIV_HE80q;_j
RRRR-RR-NRD#P0RCFO0sR
RRRRRL0Hos5CCI0H8EIq*HE800R-48MFI05FRI0H8E4q-2H*I800E2=R<RmRBh1e_ap7_mBtQ_Be a5m)j4,R2R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR&RRRo#HMR4
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR&ARq58IH0*EAI0H8E4q-RI8FMR0FI0H8E5A*I0H8E4q-2R2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR&
RqRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRB&Rm_he1_a7pQmtB _eB)am5Rj,I0H8E4q-2
;
RRRRRFRVsFDFbVd:F[sRRRHM4FR0Rb8C0oERCsMCN
0CRRRRRRRRR:l4RDRVF_FsNC88sR
RRRRRRRRRRCRoMHCsONRlb
R5RRRRRRRRRRRRRRRRRRRRR8IH0hEQR>R=ROPCD5Hl[-2RROPCD5Hl[2-4,R
RRRRRRRRRRRRRRRRRRIRRHE80mRza=P>RCHODl+5[4-2RROPCD5Hl[
2,RRRRRRRRRRRRRRRRRRRRRlMkLRCsR>R=RlMkL#Cs54[-2R
RRRRRRRRRR
R2RRRRRRRRRRRRb0FsRblNRR5
RRRRRRRRRRRRRRRRRRRRQkMb0RRRRR=>L0Hos5CCPDCOH[l52R-48MFI0PFRCHODl-5[4,22
RRRRRRRRRRRRRRRRRRRRkRm00bkR=RR>HRLoC0sCC5POlDH54[+2R-48MFI0PFRCHODl25[2R
RRRRRRRRRR;R2
RRRRCRRMR8RoCCMsCN0RsVFDbFFdR;
RMRC8CRoMNCs0HCRVF_M0C	Cb8_N8aCss;CC
R
RRFbs80kORR<=L0Hos5CCPDCOH8l5CEb0+-42.FR8IFM0ROPCD5Hl80CbE42+2
;R
8CMRONsE
4;
LDHs$NsRCHCCk;
#HCRC3CC#_08DHFoO4_4nNc3D
D;kR#CHCCC38#0_oDFHNO_sEH03DND;#
kCCRHC#C30D8_FOoH_o#HM3C8N;DD
H
DLssN$sRFO;Nd
Ck#ROFsNFd3sOONF3lbN;DD
H
DLssN$$R#MHbDV
$;kR#C#b$MD$HV30N0skHL03C#N;DD
M
C0$H0RN#lDkDvDH0R#R
RRMoCCOsH5R
RRRRRN8IH0:ERR0HMCsoCRR:=gR;
RRRRRHLI8R0E:MRH0CCos=R:R
g;RRRRRHRI8R0ERH:RMo0CC:sR=UR4
RRR2R;
RFRbs50R
RRRRqRRRRRR:MRHR0R#8F_Do_HOP0COFNs5I0H8ER-48MFI0jFR2R;
RRRRRRARRRR:HRMR#_08DHFoOC_POs0F5HLI8-0E4FR8IFM0R;j2
RRRRuRR)Rm7:kRF00R#8F_Do_HOP0COFIs5HE80-84RF0IMF2Rj
RRRR-RR-RRA*
RqR2RR;R
RR0N0skHL0\CR3lsCF_PCMIF_N\sMRH:RMo0CC
s;RNRR0H0sLCk0Rs\3N\M	RH:RMo0CC
s;CRM8#DlNDDvk0
;
NEsOHO0C0CksRONsEF4RVlR#NvDDkRD0H
#
RVRRk0MOHRFM#5kbI0H8ERN,I0H8E:LRR0HMCsoC2CRs0MksR0HMCsoCR
H#RLRRCMoH
RRRRHRRVIR5HE80NRR>I0H8ERL20MEC
RRRR0sCkRsMI0H8E
N;RRRRRDRC#RC
RsRRCs0kMHRI8L0E;R
RRRRRCRM8H
V;RCRRM#8Rk
b;
RRRVOkM0MHFRVHM58IH0,ENR8IH0REL:MRH0CCoss2RCs0kMMRH0CCos#RH
RRRLHCoMR
RRRRRH5VRI0H8E<NRR8IH02ELRC0EMR
RRCRs0MksR8IH0;EN
RRRRCRRD
#CRsRRCs0kMHRI8L0E;R
RRRRRCRM8H
V;RCRRMH8RM
V;
RRRO#FM00NMR8IH0REq:MRH0CCos=R:RVHM5HNI8,0ERHLI820E;R
RRMOF#M0N0HRI8A0ERH:RMo0CC:sR=kR#bI5NHE80,IRLHE802
;
RORRFFlbM0CMRswH#s0uFO8k0S#
SMoCCOsH5S
SS8IH0REq:MRH0CCosS;
SHSI8A0ERH:RMo0CCSs
S;S2
bSSFRs05S
SSRqR:MRHR0R#8F_Do_HOP0COFNs5I0H8ER-48MFI0jFR2S;
SRSARH:RM#RR0D8_FOoH_OPC05FsL8IH04E-RI8FMR0Fj
2;SqSSARR:FRk0#_08DHFoOC_POs0F5HLI8*0EN8IH04E-RI8FMR0FjS2
S-S-R*ARRSq
S;S2
RRRCRM8ObFlFMMC0
;
RORRFFlbM0CMR8N8CssaC
C.SCSoMHCsOS5
SHSI8q0ERH:RMo0CC
s;SISSHE80ARR:HCM0o;Cs
SSS0CsCR:RRR0HMCsoC
SSS2S;
SsbF0
R5SqSS,lRq,RRA:MRHR8#0_oDFH
O;SqSSA:RRRRHM#_08DHFoOC_POs0F5HLI8*0EN8IH04E-RI8FMR0Fj
2;SbSSskF8O:0RR0FkR8#0_oDFHPO_CFO0sI5LHE80+HNI8-0E4FR8IFM0R
j2S-SS-RRA*
RqS2SS;R
RR8CMRlOFbCFMM
0;
RRR#MHoNNDR_GNkR#:R0D8_FOoH_OPC05FsI0H8E4q-RI8FMR0Fj
2;R#RRHNoMD_RLNRkG:0R#8F_Do_HOP0COFIs5HE80AR-48MFI0jFR2R;
RHR#oDMNRRNLR:RRR8#0_oDFHPO_CFO0sI5NHE80*HLI8-0E4FR8IFM0R;j2
RRR#MHoN)DRCD#k0#:R0D8_FOoH_OPC05FsN8IH0LE+I0H8ER-48MFI0jFR2L;
CMoHRR
RRR--1bINRNqRMA8RRRHVMCCO#s#N$R
RRqHVDoNsC:sARRHV5HNI8R0E>IRLHE802CRoMNCs0RC
RRRRRsVFDbFF.V:RFHsRRRHMjFR0RHLI8-0E4CRoMNCs0RC
RRRRRRRRNs00H0LkC3R\s	NM\VRFRosC#:qRRLDNCHDR#;Rj
RRRRRRRR0RN0LsHkR0C\C3slCFP__MFIMNs\VRFRosC#:qRRLDNCHDR#;R4
RRRRRRRR0RN0LsHkR0C\N3sMR	\FsVRCAo#RD:RNDLCRRH#jR;
RRRRRRRRNs00H0LkC3R\sFClPMC_FN_IsRM\FsVRCAo#RD:RNDLCRRH#4R;
RRRRRoLCHRM
RRRRRosC#Rq:bCHbL
kVRRRRRFRbsl0RN
b5RRRRRRRRR=QR>5RAH
2,RRRRRRRRR=mR>_RNN5kGHR2
RRRRR
2;RRRRRCRso:#ARbbHCVLk
RRRRbRRFRs0l5Nb
RRRRRRRRRRQ=q>R5,H2
RRRRRRRRRRm=L>R_GNk5
H2RRRRR;R2
RRRRCRRMo8RCsMCNR0CVDFsF.Fb;R
RRRRRVDFsF4Fb:FRVsRRHHLMRI0H8EFR0RHNI8-0E4CRoMNCs0RC
RRRRRRRRNs00H0LkC3R\s	NM\VRFRosC#:ARRLDNCHDR#;Rj
RRRRRRRR0RN0LsHkR0C\C3slCFP__MFIMNs\VRFRosC#:ARRLDNCHDR#;R4
RRRRLRRCMoH
RRRRsRRCAo#:HRbbkCLVR
RRRRRb0FsRblN5R
RRRRRRQRRRR=>q25H,R
RRRRRRmRRRR=>Lk_NG25H
RRRR2RR;R
RRRRRCRM8oCCMsCN0RsVFDbFF4R;
RMRC8CRoMNCs0HCRVNqDssoCA
;
RHRRVlq#NCDDsRA:H5VRN8IH0<ER=IRLHE802CRoMNCs0RC
RRRRRsVFDbFFNV:RFHsRRRHMjFR0RHNI8-0E4CRoMNCs0RC
RRRRRRRRNs00H0LkC3R\s	NM\VRFRosC#:BRRLDNCHDR#;Rj
RRRRRRRR0RN0LsHkR0C\C3slCFP__MFIMNs\VRFRosC#:BRRLDNCHDR#;R4
RRRRRRRR0RN0LsHkR0C\N3sMR	\FsVRC1o#RD:RNDLCRRH#jR;
RRRRRRRRNs00H0LkC3R\sFClPMC_FN_IsRM\FsVRC1o#RD:RNDLCRRH#4R;
RRRRRoLCHRM
RRRRRosC#RB:bCHbL
kVRRRRRFRbsl0RN
b5RRRRRRRRR=QR>5RqH
2,RRRRRRRRR=mR>_RNN5kGHR2
RRRRR
2;RRRRRCRso:#1RbbHCVLk
RRRRbRRFRs0l5Nb
RRRRRRRRRRQ=A>R5,H2
RRRRRRRRRRm=L>R_GNk5
H2RRRRR;R2
RRRRCRRMo8RCsMCNR0CVDFsFNFb;R
RRRRRVDFsFLFb:FRVsRRHHNMRI0H8EFR0RHLI8-0E4CRoMNCs0RC
RRRRRRRRNs00H0LkC3R\s	NM\VRFRosC#:7RRLDNCHDR#;Rj
RRRRRRRR0RN0LsHkR0C\C3slCFP__MFIMNs\VRFRosC#:7RRLDNCHDR#;R4
RRRRLRRCMoH
RRRRsRRC7o#:HRbbkCLVR
RRRRRb0FsRblN5R
RRRRRRQRRRR=>A25H,R
RRRRRRmRRRR=>Lk_NG25H
RRRR2RR;R
RRRRRCRM8oCCMsCN0RsVFDbFFLR;
RMRC8CRoMNCs0HCRVlq#NCDDs
A;
RRRw#Hs0C10bw:RH0s#u8sFk#O0
RRRoCCMsRHOlRNb5R
RRRRRI0H8E=qR>HRI8q0E,R
RRRRRI0H8E=AR>HRI8A0E
RRR2R
RRsbF0NRlb
R5RRRRRRRq=N>R_GNk,R
RRRRRA>R=RNL_k
G,RRRRRARqRR=>NRL
R;R2
R
RR8q8CssaC:CRR8N8CssaC
C.RoRRCsMCHlORN5bR
RRRRIRRHE80q>R=R8IH0,Eq
RRRRIRRHE80A>R=R8IH0,EA
RRRR0RRsRCCR>R=RRjRRRRRRR--4VRHR8N8CNsRVs0CRC0ERDlk0DHbH,CsRCjRD
#CR2RR
RRRb0FsRblNRR5
RRRRRRql=N>R_GNk5,j2
RRRRqRRR>R=RNN_kIG5HE80q2-4,R
RRRRRA=RR>_RLN5kGI0H8E4A-2R,
RRRRRRqA=N>RLR,
RRRRRFbs80kORR=>)kC#DR0
R;R2
R
RR_HVIRF:H5VRI0H8E=R<R8IH0REq+HRI8A0E2CRoMNCs0RC
RRRRRmu)7=R<R#)Ck5D0I0H8ER-48MFI0jFR2R;
RMRC8CRoMNCs0HCRVF_I;R
RR_HVIR4:H5VRI0H8ERR>I0H8E+qRR8IH02EARMoCC0sNCR
RRRRRu7)m58IH0+EqI0H8E4A-RI8FMR0Fj<2R=CR)#0kD58IH0+EqI0H8E4A-RI8FMR0Fj
2;RRRRRFRVsF_DFIb_:FRVsRRHHIMRHE80qH+I8A0ERR0FI0H8ER-4oCCMsCN0
RRRRRRRR)RumH752=R<R#)Ck5D0I0H8EIq+HE80A2-4;R
RRRRRCRM8oCCMsCN0RsVF_FDFb;_I
RRRCRM8oCCMsCN0R_HVI
4;CRM8NEsO4
;
-*-R*************************************************************R**R
---e-R.mApBqi5,,RARmu)7-2
--
-RHNI8R0E-HRI8R0EFqVRRbHMk-0
-IRLHE80RI-RHE80RRFVAMRHb
k0-
-R-u-R)Rm7-ERaCkRVDbDRskF8O50RN8IH0+ERRHLI8R0EICH82sRVFLlRD	FORDlk0DHbH#Cs3-R
--R
-*R**************************************************************R*R-
-
DsHLNRs$HCCC;#
kCCRHC#C30D8_FOoH_n44cD3NDk;
#HCRC3CC#_08DHFoOs_NH30EN;DD
Ck#RCHCC03#8F_Do_HOkHM#o8MC3DND;D

HNLssF$RsdON;#
kCsRFO3NdFNsOObFl3DND;C

M00H$.ReABpmi#RH
CSoMHCsO
R5SNSSI0H8ERR:HCM0o;Cs
SSSL8IH0:ERR0HMCsoC;S
SSCMC8H_bbkCLV:#RR0HMCsoC2S;
b0FsRS5
SRqRRRR:HRMR#_08DHFoOC_POs0F5HNI8-0E4FR8IFM0R;j2
ASSRRRR:MRHR0R#8F_Do_HOP0COFLs5I0H8ER-48MFI0jFR2S;
Smu)7RR:FRk0#_08DHFoOC_POs0F5HNI8+0EL8IH04E-RI8FMR0Fj;22
0SN0LsHkR0C\N3sMR	\:MRH0CCosS;
Ns00H0LkC3R\sFClPMC_FN_IsRM\:MRH0CCosS;
Ns00H0LkC3R\LHCoMs_0CRC\:MRH0CCosS;
Ns00H0LkC3R\HCM0sDMN_#HM00NMHCN08:\RR0HMCsoC;M
C8.ReABpmi
;
NEsOHO0C0CksRFLDOR	#FeVR.mApBHiR#S

-q-RRGlNHllkRMVkOF0HMCRMC88CRCIEMIRNHE80RRH#MRF0CNJkDFR0RHLI8
0ESR--bbksF:#CRMVH8ER0CJR#kCNsRsNsNI$RHE80RFVslER0CMRHbRk0LRk##CHx#R
RRMVkOF0HM$RllRNG5DPNk,CNRDPNkRCL:MRH0CCosS2
S0sCkRsMHCM0oRCsHS#
LHCoM-RR-$Rll
NGSVSHRDPNkRCN>NRPDLkCRC0EMS
SS0sCkRsMPkNDC
N;SDSC#SC
SCSs0MksRDPNk;CL
CSSMH8RVS;
CRM8lN$lG
;
SR--bbksF:#CRDBNONkD00CREHCRMG8CRRHM0RECu8sFkRO0qNss$VRFRC0ER0CMsS$
-0-RERN08CC0sMlHC0#RE#CRHRoMLRH0VRFs0RECOsksCRM0s3FIRR
RRMVkOF0HMHR1oDMAFRO	5R
RRRRRO#FM00NMR8IHNI,RH,8LRGH8RH:RMo0CC
s2SCSs0MksR0HMCsoCR
H#SoLCHRMR-1-RHAoMD	FO
HSSVIR5H-8N4H2-8<GRR8IHLER0CSM
SCSs0MksRI55H+8L452*INH8--42H28G;S
SCCD#
SSSskC0s5MRILH8*H5I8HL+8-G24
2;SMSC8VRH;C
SM18RHAoMD	FO;R

RFROlMbFCRM0vazp44UXUv_ 
RRRRbRRFRs05S
Sq,4(Rnq4,4Rq6q,R4Rc,q,4dR.q4,4Rq4q,R4Rj,qRgRRRRRR:RRRRHM#_08DHFoO
R;SUSq,(Rq,nRq,6Rq,cRq,dRq,.Rq,4Rq,jRqSSSSR:RRRRHM#_08DHFoO
R;S4SA(A,R4Rn,A,46RcA4,4RAdA,R4R.,A,44RjA4,gRARRRRRRRRRH:RM0R#8F_DoRHO;S
SARU,AR(,ARn,AR6,ARc,ARd,AR.,AR4,ASjSSRSRRH:RM0R#8F_DoRHO;S

RRRRu,d6Rcud,dRudu,RdR.,u,d4Rjud,.Rugu,R.RU,uR.(RRRRR:RRR0FkR8#0_oDFH;OR
uSS.Rn,u,.6Rcu.,.Rudu,R.R.,u,.4Rju.,4Rugu,R4SUSR:RRR0FkR8#0_oDFH;OR
uSS4R(,u,4nR6u4,4Rucu,R4Rd,u,4.R4u4,4Ruju,RgRRRRRRRRRR:FRk0#_08DHFoO
R;SUSu,(Ru,nRu,6Ru,cRu,dRu,.Ru,4Ru,jRuSSSSR:RRR0FkR8#0_oDFH
ORS;S2
MSC8FROlMbFC;M0
R
RRMOF#M0N0zRWvRRRRH:RMo0CC:sR=(R4;-R-R8IH0FERVsRFOkNdMo#HMRC8LODF	kRlDb0HDsHC
RRRO#FM00NMRvW1RRRR:MRH0CCos=R:R;4URR--I0H8EVRFROFsNHd#o8MCRFLDOl	RkHD0bCDHsR

RFROMN#0MZ0R 4)m(RR:#_08DHFoOC_POs0FRR:="jjjjjjjjjjjjjjjj;j"
O
SF0M#NRM0INH8R:RRR0HMCsoCRR:=5I5NHE80+vWz-/.2W2zv;-RR-HR#oLMRHH0R#sR8FCbb8R
RRMOF#M0N0HRI8RLRRH:RMo0CC:sR=5R5L8IH0WE+z.v-2z/WvR2;RR--#MHoR0LHRRH#8bsFb
C8RORRF0M#NRM0I8bsR:RRR0HMCsoCRR:=INH8RI+RH;8LR-R-R8IH0FERVsRbFO8k0O
SF0M#NRM0IsNsR:RRR0HMCsoCRR:=INH8RI*RH;8LR-R-R8IH0FERVNRusN0HDsRuFO8k0sRNs
N$RORRF0M#NRM0IGlNR:RRR0HMCsoCRR:=lN$lGH5I8RN,ILH82
;
SR--aRECHkMb0N#Rs#CRb0DHR0HMF(R4-0LHRkOEM,	#RC0EMNRCOOERE	kMRRH##MHoR0CGCCM88R
RRb0$C0Rq$RbCHN#Rs$sNRR5j0IFRH-8N4F2RV0R#8F_Do_HOP0COFRs5RvW1-84RF0IMF2Rj;R
RRb0$C0RA$RbCHN#Rs$sNRR5j0IFRH-8L4F2RV0R#8F_Do_HOP0COFRs5RvW1-84RF0IMF2Rj;

RSR--0RECClDCC#M0RRFV0RECu0NsHRND1Rkl)#FIRCNsR-4(L#H0R8IHCR
RRb0$C0R1$RbCHN#Rs$sNRR5j0IFRb-s84F2RV0R#8F_Do_HOP0COFRs5RvWz-84RF0IMF2Rj;S

-0-REbCRNHs0NbDRskF8OR0#NRsCdLn-HR0#ICH8
RRR0C$bR$u0bHCR#sRNsRN$50jRFNRIs4s-2VRFR8#0_oDFHPO_CFO0s*5.W-1v4FR8IFM0R;j2
-
S-ERaCMRHb#k0RRHMNHRI8NNRs$sNRRFV4LU-HO0RE	kM##
SHNoMDNRqs$sNRRRR:0Rq$;bC
HS#oDMNRsANsRN$R:RRR$A0b
C;
-S-RC0ERsuN0DHNRFus80kORsNsNN$R#RRNIsNsRsNsNF$RVnRd-0LHRkOEM
	#R#RRHNoMDLRukRVRRRRR:0Ru$;bC
RRR#MHoNuDRsqF8s$sNRu:R0C$b;

SLHCoM-RR-DRLF#O	
-
S-ERaCR#C0RIFbOsFCC###ERONCMoRC0ERsPNHDNLCHRI8R0EHkMb0H#RMR0FVCHG8HRI8R0EHkMb0
#3SR--aRECI0H8EVRFRC0ERbHMkR0#NRsCHWMR1ovRsbFk#FRVsFRL0RE3RI]FCsPC,ER0CUR4-0LH
-S-RFoskRb#CENORMOF0MNHRR4(L#H0RFVslER0CsRFHMoHNRD,CCGObV0RF0sRElCRF
#0SR--#MHoHOVHNRM0oksFbER0NN0RDR#FERN#0REC#MHoR0LHRRFV0RECFosHHDMN3R
RR#sCH_xCNb:RsCFO#5#RqS2
PHNsNCLDR0 GqDeNS:RRR8#0_oDFHPO_CFO0s15WvR-48MFI0jFR2S;
LHCoM-RR-sRbF#OC#CRs#CHx_RN
RRRRRsVFRGH8RRHMjFR0RvW1-D4RF
FbSHSSVIR5H-8N4W2*zHv+8NG<I0H8EER0CRMR-O-RFRb$FosHHDMNR0LH#S
SSGS 0NqeD85HG:2R=5Rq5H5I84N-2z*WvH2+8;G2
SSSCCD#RRSS-#-RHRoMCCG0MS8
S SSGe0qNHD58RG2:q=R5Dq'C2V0;S
SS8CMR;HV
CSSMD8RF;FbR-R-RGH8
qSSNNss$H5I84N-2=R<R0 GqDeN;S
S-8-RFFRM0HR#oCMRGM0C81RpAsRoF#kb
VSSFHsR8HGRMRRj0IFRH-8N.FRDFSb
SNSqs$sN5GH82=R<R''jRq&R5vWz*85HG2+4-84RF0IMFzRWv8*HG
2;RRRRRMRC8FRDF
b;S8CMRFbsO#C#R#sCH_xCN
;
RsRRCx#HC:_LRFbsO#C#R25A
NSPsLHND CRGe0ANRDSR#:R0D8_FOoH_OPC05FsW-1v4FR8IFM0R;j2
RRRLHCoM-RR-sRbF#OC#CRs#CHx_RL
RRRRRsVFRGH8RRHMjFR0RvW1-D4RF
FbSHSSVIR5H-8L4W2*zHv+8LG<I0H8EER0CRMR-O-RFRb$FosHHDMNR0LH#S
SSGS 0NAeD85HG:2R=5RA5H5I84L-2z*WvH2+8;G2
SSSCCD#RRSS-#-RHRoMCCG0MS8
S SSGe0ANHD58RG2:A=R5DA'C2V0;S
SS8CMR;HV
CSSMD8RF;FbR-R-RGH8
ASSNNss$H5I84L-2=R<R0 GADeN;S
S-8-RFFRM0HR#oCMRGM0C81RpAsRoF#kb
RRRRVRRFHsR8HGRMRRj0IFRH-8L.FRDFSb
SNSAs$sN5GH82=R<R''jRA&R5vWz*85HG2+4-84RF0IMFzRWv8*HG
2;SMSC8FRDFRb;RR--H
8GRCRRMb8RsCFO#s#RCx#HC;_L
-
S-CRoMNCs00CREuCRNHs0NuDRskF8ON0Rs$sNRRL$l0kDH$bDHRMo0REC4LU-HO0RE	kM#VRF
-S-RC0ERbHMkR0#0VFRFRsldLn-Hu0RNHs0NuDRskF8O30#R
R
SMoCl0kDNV:RFNsRGMRHR0jRFHRI84N-RMoCC0sNCS
SolCMkLD0:FRVsGRLRRHMjFR0R8IHLR-4oCCMsCN0
SSSNs00H0LkC3R\HCM0sDMN_#HM00NMHCN08F\RVkRlDG0GRD:RNDLCRRH#4S;
SoLCHSM
SkSlDG0GRv:Rz4paUUX4_
 vRRRRRFRbsl0RN5bR
RRRRRRRR4Rq(>R=RsqNs5N$N5G24,(2
RRRRRRRR4Rqn>R=RsqNs5N$N5G24,n2
RRRRRRRR4Rq6>R=RsqNs5N$N5G24,62
RRRRRRRR4Rqc>R=RsqNs5N$N5G24,c2
RRRRRRRR4Rqd>R=RsqNs5N$N5G24,d2
RRRRRRRR4Rq.>R=RsqNs5N$N5G24,.2
RRRRRRRR4Rq4>R=RsqNs5N$N5G24,42
RRRRRRRR4Rqj>R=RsqNs5N$N5G24,j2
RRRRRRRRgRqRR=>qsNsNN$5Gg252R,
RRRRRRRRq=UR>NRqs$sN52NG5,U2
RRRRRRRR(RqRR=>qsNsNN$5G(252R,
RRRRRRRRq=nR>NRqs$sN52NG5,n2
RRRRRRRR6RqRR=>qsNsNN$5G6252R,
RRRRRRRRq=cR>NRqs$sN52NG5,c2
RRRRRRRRdRqRR=>qsNsNN$5Gd252R,
RRRRRRRRq=.R>NRqs$sN52NG5,.2
RRRRRRRR4RqRR=>qsNsNN$5G4252R,
RRRRRRRRq=jR>NRqs$sN52NG5,j2
RRRRRRRR4RA(>R=RsANs5N$L5G24,(2
RRRRRRRR4RAn>R=RsANs5N$L5G24,n2
RRRRRRRR4RA6>R=RsANs5N$L5G24,62
RRRRRRRR4RAc>R=RsANs5N$L5G24,c2
RRRRRRRR4RAd>R=RsANs5N$L5G24,d2
RRRRRRRR4RA.>R=RsANs5N$L5G24,.2
RRRRRRRR4RA4>R=RsANs5N$L5G24,42
RRRRRRRR4RAj>R=RsANs5N$L5G24,j2
RRRRRRRRgRARR=>AsNsNL$5Gg252R,
RRRRRRRRA=UR>NRAs$sN52LG5,U2
RRRRRRRR(RARR=>AsNsNL$5G(252R,
RRRRRRRRA=nR>NRAs$sN52LG5,n2
RRRRRRRR6RARR=>AsNsNL$5G6252R,
RRRRRRRRA=cR>NRAs$sN52LG5,c2
RRRRRRRRdRARR=>AsNsNL$5Gd252R,
RRRRRRRRA=.R>NRAs$sN52LG5,.2
RRRRRRRR4RARR=>AsNsNL$5G4252R,
RRRRRRRRA=jR>NRAs$sN52LG5,j2
RRRRRRRRdRu6>R=RkuLVN55GH*I8+L2L5G2d,62
RRRRRRRRdRuc>R=RkuLVN55GH*I8+L2L5G2d,c2
RRRRRRRRdRud>R=RkuLVN55GH*I8+L2L5G2d,d2
RRRRRRRRdRu.>R=RkuLVN55GH*I8+L2L5G2d,.2
RRRRRRRRdRu4>R=RkuLVN55GH*I8+L2L5G2d,42
RRRRRRRRdRuj>R=RkuLVN55GH*I8+L2L5G2d,j2
RRRRRRRR.Rug>R=RkuLVN55GH*I8+L2L5G2.,g2
RRRRRRRR.RuU>R=RkuLVN55GH*I8+L2L5G2.,U2
RRRRRRRR.Ru(>R=RkuLVN55GH*I8+L2L5G2.,(2
RRRRRRRR.Run>R=RkuLVN55GH*I8+L2L5G2.,n2
RRRRRRRR.Ru6>R=RkuLVN55GH*I8+L2L5G2.,62
RRRRRRRR.Ruc>R=RkuLVN55GH*I8+L2L5G2.,c2
RRRRRRRR.Rud>R=RkuLVN55GH*I8+L2L5G2.,d2
RRRRRRRR.Ru.>R=RkuLVN55GH*I8+L2L5G2.,.2
RRRRRRRR.Ru4>R=RkuLVN55GH*I8+L2L5G2.,42
RRRRRRRR.Ruj>R=RkuLVN55GH*I8+L2L5G2.,j2
RRRRRRRR4Rug>R=RkuLVN55GH*I8+L2L5G24,g2
RRRRRRRR4RuU>R=RkuLVN55GH*I8+L2L5G24,U2
RRRRRRRR4Ru(>R=RkuLVN55GH*I8+L2L5G24,(2
RRRRRRRR4Run>R=RkuLVN55GH*I8+L2L5G24,n2
RRRRRRRR4Ru6>R=RkuLVN55GH*I8+L2L5G24,62
RRRRRRRR4Ruc>R=RkuLVN55GH*I8+L2L5G24,c2
RRRRRRRR4Rud>R=RkuLVN55GH*I8+L2L5G24,d2
RRRRRRRR4Ru.>R=RkuLVN55GH*I8+L2L5G24,.2
RRRRRRRR4Ru4>R=RkuLVN55GH*I8+L2L5G24,42
RRRRRRRR4Ruj>R=RkuLVN55GH*I8+L2L5G24,j2
RRRRRRRRgRuRR=>uVLk5G5N*8IHLL2+Gg252R,
RRRRRRRRu=UR>LRuk5V5NIG*H28L+2LG5,U2
RRRRRRRR(RuRR=>uVLk5G5N*8IHLL2+G(252R,
RRRRRRRRu=nR>LRuk5V5NIG*H28L+2LG5,n2
RRRRRRRR6RuRR=>uVLk5G5N*8IHLL2+G6252R,
RRRRRRRRu=cR>LRuk5V5NIG*H28L+2LG5,c2
RRRRRRRRdRuRR=>uVLk5G5N*8IHLL2+Gd252R,
RRRRRRRRu=.R>LRuk5V5NIG*H28L+2LG5,.2
RRRRRRRR4RuRR=>uVLk5G5N*8IHLL2+G4252R,
RRRRRRRRu=jR>LRuk5V5NIG*H28L+2LG5
j2S;S2
S
SS_HVbLHb4H:RVMR5C_C8bCHbL#kVR4=R2CRoMNCs0SC
SLSSkbVbHV:RFHsRRRHMjFR0RW.*14v-RMoCC0sNCS
SSNSS0H0sLCk0Rs\3N\M	RRFVs#CoRD:RNDLCRRH#4S;
SSSSNs00H0LkC3R\LHCoMs_0CRC\FsVRCRo#:NRDLRCDH4#R;S
SSNSS0H0sLCk0Rs\3CPlFCF_M_sINMF\RVCRso:#RRLDNCHDR#;R4
SSSSoLCH
MRSSSSSosC#R:RbCHbL
kVSSSSSsbF0NRlbS5
SSSSSRSQ=u>RL5kV5*NGILH82G+L225H,S
SSSSSS=mR>sRuFs8qs5N$5*NGILH82G+L225H2S;
SCSSMo8RCsMCNR0CLbkVb
H;SCSSMo8RCsMCNR0CHbV_H4bL;S
SS_HVbLHbjH:RVMR5C_C8bCHbL#kVRj=R2CRoMNCs0SC
SuSSsqF8s$sN5G5N*8IHLL2+G<2R=LRuk5V5NIG*H28L+2LG;S
SS8CMRMoCC0sNCVRH_bbHL
j;SMSC8CRoMNCs0oCRCkMlD;0L
MSC8CRoMNCs0oCRCkMlD;0N
-
S-NRa	0CREuCRNHs0NuDRskF8ON0Rs$sNR8NMRHLkD08RENCR8s8CRC0sCR3RqkRsMMMHokR#l-
S-#RHRHHM0HNDx,C8RC0EM0RFERCss#FIRRFV0RECb0NsHRNDb8sFkRO0NRsCNC888S3
-w-RFCsRGbNlDRC,HqVRRRH#6LU-HR0#ICH8R8NMRHAR#cR.-0LH#HRI8RC,0MECRVqRHR0#HcMR
-S-R-4(LRH0OMEk	N#RMA8RR0VH#MRHR4.R(H-L0EROk#M	3aRRENCRs$sNRDIHDMRHO8DkC*Rc.S=
-U-RRDlk0DHbH#CsRsVFloHMRdURnH-L0NRusN0HDsRuFO8k0R#3RCaERDVkDsRbFO8k0HRIDLDRCSR
-c-R+n.=R-4(LRH0OMEk	I#RH38CRERaCkR)Ml1kRRH#H0MHHHNDxRC80
F:SR--R1RRH oMGR0,RHR1oGM 0R,RR5uu42,4ERH,u4u5,D42Fu,Ru,5jjH2E,uRu5jj,2
DFSR--aMECREF0CssRFRI#NRsCVlFsCL8RN8#CRRFM0RECI0H8EVRFRHqRM(R4-0LHRkOEMR	#N
M8SR--0RECI0H8EVRFRHARM(R4-0LHRkOEM3	#RFRwsER0CGRCNDlbCS:
-a-RE'CRqD'RFRFb504RF2Rd
-S-RRRR1MHo ,G0RuRRu,5.4H2E,uRu54.,2,DFR5uu42,jERH,u4u5,Dj2Fj,R'S#
-R-RRuRu54d,2,EHR5uud2,4DRF,u.u5,Ej2Hu,Ru,5.jF2D,'Rj#R,RRRRRR#j'
-S-RRRR1MHo ,G0RuRRu,5djH2E,uRu5jd,2,DFR#j',RRRRRRRj,'#RRRRRjRR'S#
-a-RE'CRAD'RFRFb504RF2R4
-S-RRRR1MHo ,G0R1RRH oMGR0,RHR1oGM 0R,RR5uuj2,4ERH,uju5,D42Fj,R'S#
-w-RFNsRRslFCER0FksFoCERGNbDMHN0FRM,#RCC0RECe0HsCQG-QDRAFRO	v0kDHHbDCSs
-#-RbHCOVNHO0MHF3
R
RNRR8s8bFR8:bOsFCR##5Fus8sqsN
$2SNSPsLHND)CRkkM1lRRRR#:R0D8_FOoH_OPC05FsI8bs*vWz+84RF0IMF2RjRR:=5EF0CRs#='>Rj;'2
RRRRPRRNNsHLRDC1)klFCIeORR:#_08DHFoOC_POs0F5sIb8z*WvR+48MFI0jFR2R;
RRRRRsPNHDNLCkR1lI)FRRRR:0R1$;bC
RRRRPRRNNsHLRDCNGH8RRRRRRR:HCM0o;Cs
RRRRPRRNNsHLRDCLGH8RRRRRRR:HCM0o;Cs
RRRRPRRNNsHLRDC[RRRRRRRRRR:HCM0o;Cs
RRRRPRRNNsHLRDC	RRRRRRRRRR:HCM0o;Cs
CSLoRHMRR--bOsFCR##Nb88s
F8S-S-RHQM0DHNHRxC0RECsMkMHRMo#Rkl5M)k12kl
RRRRVRRFNsRGMRHR0jRFlRIN4G-RFDFbS
SS8LHG=R:R;NG
SSS[RRRRR:=.G*N;S
SSR	RR=R:R+[RR
4;SHSSVGRNRI>RH-8N4sRFR8LHGRR>ILH8-04RE
CMSSSSH[VRRI<RbRs80MECRSRSRR--#MHoR0CGC
M8SSSSSl1k)5FI[:2R=FR50sEC#>R=RFus8sqsN1$5HAoMD	FO58IHNH,I8jL,2.25*vW1-2.2;S
SSMSC8VRH;S
SSVSHR<	RRsIb8ER0CRMRS-SR-HR#oCMRGM0C8S
SS1SSkFl)I25	RR:=5EF0CRs#=u>RsqF8s$sN5o1HMFADOI	5H,8NILH8,2j25W.*1.v-2
2;SSSSCRM8H
V;SCSSD
#CSSSS1)klF[I52=R:RFus8sqsNN$5GH*I8LL+H28G5WRRz4v-RI8FMR0FR2Rj;R
RRRRRRRRRRVRHR<	RRsIb8ER0CSM
SSSS1)klF	I52=R:RFus8sqsNN$5GH*I8LL+H28G5W.*z4v-RI8FMR0FW2zv;S
SSMSC8VRH;S
SS8CMR;HV
SSS-O-RFCMPs00RENCRs$sNRRFVOMEk	H#RMR0FNNMRs$sNRRFVL#H0
SSSVRFsHRLGHjMRRR0FI8bs-D4RF
FbSSSSVRFsDHGRMRRj0WFRz4v-RFDFbS
SS)SSkkM1lL5HGz*WvG+D2=R:Rl1k)5FIH2LG52DG;S
SSMSC8FRDFRb;RR--DSG
SMSC8FRDFRb;RR--H
LGS-SS-MRHHN0HDCHxRC0ERo#HMHRL0S#
SkS)Ml1k5sIb8z*WvR+48MFI0IFRb*s8W2zvRR:=5EF0CRs#=u>RsqF8s$sN5o1HMFADOI	5H,8NILH8,2j25W.*1.v-2
2;SMSC8FRDFRb;RR--NSG
SR--pbFFRRFM0RECqMRH8
CGSFSVs8RHGMRHR04RFHRI84N-RFDFbR
RRRRRRVRRFNsRGMRHR0jRFlRIN4G-RFDFbS
SSHSL8:GR=GRNRH-R8
G;SSSS[RRRRR:=N+GRR8LHGS;
S	SSRRRR:[=RR4+R;S
SSVSHRRNG>HRI84N-RRFsLGH8RI>RH-8L4ER0CRM
RRRRRRRRRRRRRVRHR<[RRsIb8ER0CRMRS-SR-HR#oCMRGM0C8S
SSSSS1)klF[I52=R:R05FE#CsRR=>5Fus8sqsN1$5HAoMD	FO58IHNH,I8HL,82G25W.*1.v-2;22
SSSSMSC8VRH;S
SSHSSVRR	<bRIs08RERCMRRSS-#-RHRoMCCG0MS8
SSSSSl1k)5FI	:2R=FR50sEC#>R=Rs5uFs8qs5N$1MHoAODF	H5I8IN,H,8LH28G2*5.W-1v.222;S
SSCSSMH8RVS;
SCSSDV#HR8LHGRR<jER0CSM
SSSSH[VRRj<RRC0EMSRRS-SR-8RN[0k#RC0ER8HMO#HCR8lFkRDFIGlN
SSSS[SSRR:=[RR+.l*IN
G;RRRRRRRRRRRRRCRRMH8RVR;
RRRRRRRRRRRRRVRHR<	RR0jRE
CMSSSSSRS	:	=RR.+R*NIlGS;
SSSSCRM8H
V;SSSSSRHV[RR<N0GRE
CMSSSSSkS1lI)F5R[2:Z=R 4)m(S;
SSSSCHD#VRR[<bRIs08RERCMRRSS-#-RHRoMCCG0MS8
SSSSSl1k)5FI[:2R=FR50sEC#>R=Rs5uFs8qs5N$1MHoAODF	H5I8IN,H,8LH28G2*5.W-1v.222;S
SSCSSMH8RVS;
SSSS-F-R0sECICH#,ER0CMRH8RCGHM#RFH0RMER0CkR1lI)F,FR8R0MFEoHM
SSSSVSHR<	R=GRNRC0EMS
SSSSS1)klF	I52=R:R)Z m;4(
RRRRRRRRRRRRRRRCHD#VRR	<bRIs08RERCMRRSS-#-RHRoMCCG0MS8
SSSSSl1k)5FI	:2R=FR50sEC#>R=Rs5uFs8qs5N$1MHoAODF	H5I8IN,H,8LH28G2*5.W-1v.222;S
SS-SS-0RFEICsH,#CRC0ER8HMCHGR#FRM0MRHRC0ERl1k),FIRR8FMEF0H
MoSSSSS8CMR;HV
SSSS#CDCSRRSSSSS-SR-FRMsDlNRFbs80kORs0ClS
SS1SSkFl)I25[RR:=u8sFqNss$G5N*8IHLH+L85G2RzRWvR-48MFI0RFRR;j2
SSSSVSHR<	RRsIb8ER0CSM
SSSSSl1k)5FI	:2R=sRuFs8qs5N$NIG*H+8LLGH82*5.W-zv4FR8IFM0RvWz2S;
SSSSCRM8H
V;SSSSCRM8H
V;SCSSMD8RF;FbR-R-R
NGS-SS-FROMsPC0ER0CsRNsRN$FOVRE	kM#MRH0NFRMsRNsRN$FLVRH
0#RRRRRRRRRsVFRGHLRRHMjFR0RsIb8R-4DbFF
SSSSsVFRRDGHjMRRR0FW-zv4FRDFSb
SSSS1)klFCIeOL5HGz*WvG+D2=R:Rl1k)5FIH2LG52DG;S
SSMSC8FRDFRb;RR--DSG
SMSC8FRDFRb;RR--H
LGS-SS-CR10ER0CHR#oLMRHR0#VRFs0#EHRIsF
RRRRRRRRkR1lI)Fe5COI8bs*vWz+84RF0IMFbRIsW8*zRv2:R=R5EF0CRs#=u>RsqF8s$sN5o1HMFADOI	5H,8NILH8,GH82.25*vW1-2.2;S
SSR--qR880RECsRFI[0k#RCOsN80CRR0F0RECsMkMHRMo#
klRRRRRRRRRM)k1Rkl:)=RkkM1lRR+1)klFCIeOS;
S8CMRFDFbR;R-H-R8SG
SR--pbFFRRFM0RECAMRH8
CGSFSVsxRHGMRHR04RFHRI84L-RFDFbR
RRRRRRVRRFLsRGMRHR0jRFlRIN4G-RFDFbS
SSHSN8:GR=GRLRH-Rx
G;SSSS[RRRRR:=NGH8RL+RGS;
S	SSRRRR:[=RR4+R;S
SSVSHRRLG>HRI84L-RRFsNGH8RI>RH-8N4ER0CRM
RRRRRRRRRRRRRVRHR<[RRsIb8ER0CRMRS-SR-HR#oCMRGM0C8S
SSSSS1)klF[I52=R:R05FE#CsRR=>5Fus8sqsN1$5HAoMD	FO58IHNH,I8-L,H2xG2*5.W-1v.222;S
SSCSSMH8RVS;
SSSSH	VRRI<RbRs80MECRSRSRR--#MHoR0CGC
M8SSSSSkS1lI)F5R	2:5=RFC0Es=#R>uR5sqF8s$sN5o1HMFADOI	5H,8NILH8,x-HG522.1*Wv2-.2
2;SSSSS8CMR;HV
SSSS#CDHNVRHR8G<RRj0MEC
SSSSVSHR<[RR0jRERCMRSSSRR--Nk8[#00REHCRMH8OCl#RFD8kFlRINSG
SSSSS:[R=RR[+*R.IGlN;S
SSCSSMH8RVS;
SSSSH	VRRj<RRC0EMS
SSSSS	=R:R+	RRI.*l;NG
SSSSMSC8VRH;S
SSHSSVRR[<GRLRC0EMS
SSSSS1)klF[I52=R:R)Z m;4(
RRRRRRRRRRRRRRRCHD#VRR[<bRIs08RERCMRRSS-#-RHRoMCCG0MS8
SSSSSl1k)5FI[:2R=FR50sEC#>R=Rs5uFs8qs5N$1MHoAODF	H5I8IN,H,8L-GHx2.25*vW1-2.22S;
SSSSCRM8H
V;SSSSSRHV	=R<RRLG0MEC
SSSS1SSkFl)I25	RR:=Zm )4
(;RRRRRRRRRRRRRCRRDV#HR<	RRsIb8ER0CRMRS-SR-HR#oCMRGM0C8S
SSSSS1)klF	I52=R:R05FE#CsRR=>5Fus8sqsN1$5HAoMD	FO58IHNH,I8-L,H2xG2*5.W-1v.222;S
SSCSSMH8RVS;
SCSSD
#CSSSSSl1k)5FI[:2R=sRuFs8qs5N$NGH8*8IHLG+L2R5RW-zv4FR8IFM0RjRR2S;
SSSSH	VRRI<RbRs80MEC
SSSS1SSkFl)I25	RR:=u8sFqNss$H5N8IG*H+8LL5G2.z*WvR-48MFI0WFRz;v2
SSSSMSC8VRH;S
SSMSC8VRH;S
SS8CMRFDFbR;R-L-RGS
SSR--OPFMCRs00RECNNss$VRFRkOEMR	#HFM0RRNMNNss$VRFR0LH#R
RRRRRRVRRFHsRNHGRMRRj0IFRb-s84FRDFSb
SVSSFDsRGMRHR0jRFzRWvR-4DbFF
SSSSkS1lI)Fe5COH*NGW+zvDRG2:1=RkFl)IN5HGD25G
2;SSSSCRM8DbFF;-RR-GRD
SSSCRM8DbFF;-RR-NRHGS
SSR--1RC00REC#MHoR0LH#FRVsER0Hs#RFRI
RRRRRRRR1)klFCIeOb5IsW8*z4v+RI8FMR0FI8bs*vWz2=R:RFR50sEC#>R=RFus8sqsN1$5HAoMD	FO58IHNH,I8-L,H2xG2*5.W-1v.;22
SSS-q-R808REsCRF[IRkR#0ONsC0RC800FREsCRkHMMM#oRkRl
RRRRRRRR)1kMk:lR=kR)Ml1kR1+RkFl)IOeC;S
SCRM8DbFF;-RR-xRHGR
RRRRRu7)mRR<=)1kMkNl5I0H8EI+LHE80-84RF0IMF2Rj;C
SMb8RsCFO#N#R8s8bF
8;
8CMRFLDO;	#
-
-R****************************************************************-RR--
-R-
-R0 MHR0$7DCON0sNHRFMVRFs#MHoCl8RkHD0bCDHs-
-R-
-RHaE##RHRC0ERHlNMMRC0$H0RsVFRC0ERo#HMRC8l0kDHHbDCRs3RCaERF0IRONsECH0Os0kC-#
-CR8VCHM8CRLDRFIkR#C0RECCHM00#HCRFNLPRC,NRM8l0k#RRLCD0N#RRHM0#EHRDVHCR3Ra
EC-0-RINFRsHOE00COk#sCRCNsRC0ERoDFHPORCHs#FNMRM08RELCRD	FORsPC#MHF3-
-R-
-R****************************************************************-RR-D

HNLssH$RC;CC
Ck#RCHCC03#8F_Do_HO4c4n3DND;#
kCCRHC#C30D8_FOoH_HNs0NE3D
D;kR#CHCCC38#0_oDFHkO_Mo#HM3C8N;DD
H
DLssN$sRFO;Nd
Ck#ROFsNFd3sOONF3lbN;DD
H
DLssN$$R#MHbDV
$;kR#C#b$MD$HV30N0skHL03C#N;DD
M
C0$H0Rz1vpHaR#R
RRCRoMHCsOR5
RRRRRHRI8R0ERH:RMo0CC:sR=cR.;R
RRRRRRHNI8R0E:MRH0CCos=R:R;4.
RRRRRRRL8IH0:ERR0HMCsoCRR:=4S.
S;R2
RRRRsbF0S5
SRRqR:RRRRHM#_08DHFoOC_POs0F5HNI8R0E-84RF0IMF2Rj;S
SRRARRRR:H#MR0D8_FOoH_OPC05FsL8IH0-ER4FR8IFM0R;j2
RSSu7)mRF:Rk#0R0D8_FOoH_OPC05FsI0H8E4R-RI8FMR0FjR2
RRRRR;R2
RRRNs00H0LkC3R\s	NM\RR:HCM0o;Cs
RRRNs00H0LkC3R\lkF8DRC\:0R#soHM;R
RR0N0skHL0\CR38bFCRl\:MRH0CCosR;
R0RN0LsHkR0C\F3b8LClkR#\:0R#soHM;R
RR0N0skHL0\CR38CM_C0sC:\RR0HMCsoC;R
RR0N0skHL0\CR3oLCH0M_s\CCRH:RMo0CC
s;RNRR0H0sLCk0Rs\3CPlFCF_M_sINM:\RR0HMCsoC;M
C8vR1z;pa
-
-R****************************************************************-RR--
-R-
-RoDFHNORsHOE00COk#sCRsVFROFsN-d
--R
-*R**************************************************************R*R-
-
NEsOHO0C0CksRoDFHFORVvR1zRpaH
#
RVRRk0MOHRFMOINDHE80LOR5F0M#NRM0IRN,I:LRR0HMCsoC2CRs0MksR0HMCsoCR
H#RRRRRNRPsLHNDsCRORM0:MRH0CCosR;
RCRLo
HMRRRRRVRHRL5IRR<=IRN20MEC
RRRRRRRRORsM:0R=LRIRR;
RRRRR#CDCRR
RRRRRRRRs0OMRR:=I;NR
RRRRCRRMH8RVR;
RRRRR0sCkRsMs0OM;R
RR8CMRDONI0H8E
L;
RRRVOkM0MHFRDONI0H8E5NRO#FM00NMR,INRRIL:MRH0CCoss2RCs0kMMRH0CCos#RH
RRRRPRRNNsHLRDCs0OMRH:RMo0CC
s;RLRRCMoH
RRRRHRRVIR5L=R<R2INRC0EMR
RRRRRRsRRORM0:I=RN
R;RRRRRDRC#
CRRRRRRRRRRMsO0=R:RRIL;R
RRRRRCRM8H
V;RRRRRCRs0MksRMsO0R;
RMRC8NROD8IH0;EN
R
RRMOF#M0N0HRI8N0ERH:RMo0CC:sR=NROD8IH05ENN8IH0RE,L8IH0;E2
RRRO#FM00NMR8IH0REL:MRH0CCos=R:RDONI0H8ENL5I0H8EL,RI0H8E
2;
RRRObFlFMMC0lR#NvDDk
D0RRRRRCRoMHCsOR5
RRRRRRRRN8IH0:ERR0HMCsoCRR;
RRRRRRRRL8IH0:ERR0HMCsoCRR;
RRRRRRRRI0H8E:RRR0HMCsoC
RRRR2RR;R
RRRRRb0FsRR5
RRRRRRRRqRRRRH:RM#RR0D8_FOoH_OPC05FsN8IH04E-RI8FMR0Fj
2;RRRRRRRRRRARRRR:HRMR#_08DHFoOC_POs0F5HLI8-0E4FR8IFM0R;j2
RRRRRRRR)Rum:7RR0FkR8#0_oDFHPO_CFO0sI5RHE80-84RF0IMF2Rj
RRRR2RR;R
RR8CMRlOFbCFMM
0;
RRR#MHoNNDR_GNkRRR:#_08DHFoOC_POs0F58IH0-EN4FR8IFM0R;j2RRR
RHR#oDMNRNL_kRGR:0R#8F_Do_HOP0COFIs5HE80LR-48MFI0jFR2
;RR#RRHNoMDCR)#0kDR#:R0D8_FOoH_OPC05FsR8IH04E-RI8FMR0Fj
2;LHCoMR
RRR--p'C0#IR#NRb
RwRQ__IN#_kbIRL:H5VRN8IH0>ER=IRLHE802CRoMNCs0RC
RRRRRNN_k<GR=;RN
RRRRLRR_GNkRR<=LR;
RMRC8CRoMNCs0QCRwN_I_b#k_;IL
R
RR_QwI#L_kIb_NH:RVLR5I0H8ERR>N8IH0RE2oCCMsCN0
RRRRNRR_GNkRR<=LR;
RRRRRNL_k<GR=;RN
RRRCRM8oCCMsCN0R_QwI#L_kIb_N
;
S_HVIR4:H5VRI0H8E=LRRR42oCCMsCN0
#SSHNoMDFROlCbDl0CM,IR0FlOFbRR:#_08DHFoOC_POs0F58IH04E-RI8FMR0Fj
2;SCSLo
HMSFSVsF_DFRb:VRFsHMRHR0jRFHRI8N0E-o4RCsMCN
0CSOSSFDlbCMlC025HRR<=MRF0Nk_NG25H;SR
S8CMRMoCC0sNCFRVsF_DF
b;SOSSFDlbCMlC0H5I8-0E4<2R=FRM0_RNN5kGI0H8E4N-2S;
SIS0FlOFb=R<RlOFblDCCRM0+4R''S;
S#sCkRD0<B=Rm_he1_a7pQmtB _eB)am5Rj,I0H8EIN+HE80LI2RERCM5NL_kjG52RR='2j'
SSSS#CDCIR0FlOFbS;
SS
Su7)mRR<=skC#DI05HE80-84RF0IMF2Rj;C
SMo8RCsMCNR0CHIV_4
;
RHRRVj_I:VRHRH5I8L0ER.=R2CRoMNCs0RC
RRRRRo#HMRNDObFlDCClMR0,0OIFFRlb:0R#8F_Do_HOP0COFIs5HE80NR-48MFI0jFR2R;
RCRLo
HMRRRRRFRVsF_DFRb:VRFsHMRHR0jRFHRI8N0E-o4RCsMCN
0CRRRRRRRRRlOFblDCC5M0H<2R=FRM0_RNN5kGHR2;
RRRRCRRMo8RCsMCNR0CV_FsDbFF;R
RRRRR0OIFFRlb<O=RFDlbCMlC0RR+';4'
R
RRRRR)kC#D<0R=mRBh1e_ap7_mBtQ_Be a5m)jN,RI0H8EI+LHE802ERIC5MRLk_NG25jR'=Rj
'2RRRRRRRRRRRRCCD#RF0IObFl58IH0-EL4&2RRF0IObFl58IH0-EL4&2RRF0IObFlRCIEMLR5_GNk5R42=4R''R2
RRRRRRRRRCRRDR#CNk_NGH5I8L0E-R42&_RNN5kGI0H8E4L-2RR&Nk_NG
R;
RRRRuRR)Rm7<)=RCD#k0H5I8-0E4FR8IFM0R;j2
RRRCRM8oCCMsCN0R_HVI
j;
RRRH.V_IR4:H5VRI0H8E>LRRR.2oCCMsCN0
RRRRlRRk4D0:#RRlDNDvazp
RRRRRRRRRRRRMoCCOsHRblNRR5
RRRRRRRRRRRRRRRRRRRRN8IH0=ER>HRI8N0E,R
RRRRRRRRRRRRRRRRRRLRRI0H8E>R=R8IH0,EL
RRRRRRRRRRRRRRRRRRRRHRI8R0ERR=>I0H8ER
RRRRRRRRRR
R2RRRRRRRRRRRRb0FsRblNRR5
RRRRRRRRRRRRRRRRRRRRq>R=RNN_k
G,RRRRRRRRRRRRRRRRRRRRR=AR>_RLN,kG
RRRRRRRRRRRRRRRRRRRR)Rum=7R>)RumR7
RRRRRRRRR2RR;R
RR8CMRMoCC0sNCVRH_4.I;C

MD8RFOoH;-

-*R**************************************************************R*R---
--R
-DRLF_O	l0kDRONsECH0Os0kCV#RFFsRsdON
R--
R--****************************************************************R-R-
s
NO0EHCkO0sLCRD	FO_Dlk0VRFRz1vpHaR#S

-b-RkFsb#RC:skC0sRM#0RECMRCII0H8ENRL#RC8FCMRG#OC#HRL0L#RCoHMRCbs#0CM
RRRVOkM0MHFR#bN#8WH05ER
RRRRORRF0M#NRM0lIF8HE80RH:RMo0CC
s;RRRRRFROMN#0MF0RDH8W8R0E:MRH0CCosS2
S0sCkRsMHCM0oRCsHS#
LHCoM-RR-NRb#H#W8
0ERRRRRVRHR8lFI0H8ERR>.ER0CRMRSR--l0F#R	0NCER0HL#RsONMES
SS0sCkRsMFWD8HE80;S
SCHD#VFRl88IH0=ERR0.RE
CMSsSSCs0kMDRF88WH0.E-;S
SCHD#VFRl88IH0=ERR04RE
CMSsSSCs0kMDRF88WH04E-;S
SCHD#VFRl88IH0=ERR0jRE
CMSsSSCs0kMDRF88WH0
E;SDSC#RCRSSSSS-S-RH0E##RHRb#kCDsVk#Fk
SSSskC0sFMRDH8W8;0E
CSSMH8RVS;
CRM8b#N#W0H8E
;
SR--skC0s4MRRRHVORNMbCHbDCHMRC0ERDlk0DHbH
CsSMVkOF0HMCRMC08_FH_bbHCDMNC5I0H8EL,RI0H8ERR:HCM0o2CsR0sCkRsMHCM0oRCsHS#
LHCoMS
SH5VR5HNI8R0E>(R42MRN8LR5I0H8ERR>42(2RC0EMS
SS0sCkRsM4S;
S8CMR;HV
sSSCs0kM;Rj
MSC8CRMC08_FH_bbHCDM
C;
RRR-V-RHRM80REC#DlNDRCsI0H8EIR5HE80RRFsN8IH0
E2RVRRk0MOHRFMH5MVI0H8EN,RI0H8ERR:HCM0o2CsR0sCkRsMHCM0oRCsHR#
RCRLo
HMRRRRRVRHRH5I8R0E<IRNHE802ER0CRM
RRRRRRRRskC0sIMRHE80;R
RRRRRCCD#
RRRRRRRRCRs0MksRHNI8;0E
RRRRCRRMH8RVR;
RMRC8MRHV
;
RVRRk0MOHRFM#MHoCF8l8H5I8R0E:MRH0CCoss2RCs0kMMRH0CCos#RH
CSLoRHMRSSSSSSSSRS
RRRRRRHVI0H8Eg<4RC0EM-SR-gR4RRH#WRzv+
R.SsSSCs0kMHRI8;0ER-RR-(R4RRH#W,zvRR46HW#Rz.v-
RRRRCRRD
#CSsSSCs0kMIR5HE80--425555I0H8E6+42(/422-4*24(;S
SRMRC8VRH;
RRS8CMRo#HMlC8F
8;
RRRO#FM00NMRvWzR:RRR0HMCsoCRR:=4R(;R-SR-HRI8R0EFkVRMo#HMRC8l0kDHHbDC
s
RORRF0M#NRM0N8IHCRR:HCM0oRCs:H=RMIV5HE80,IRNHE802S;
O#FM00NMRHLI8:CRR0HMCsoCRR:=H5MVI0H8EL,RI0H8E
2;
RRRO#FM00NMRFNl8:RRR0HMCsoCRR:=#MHoCF8l8I5NH28C;R
RRMOF#M0N0lRLFR8R:MRH0CCos=R:Ro#HMlC8FL85ICH82
;
RORRF0M#NRM0N8IHRH:RMo0CC:sR=NRb#H#W850EN8lF,IRNH28C;R
RRMOF#M0N0IRLH:8RR0HMCsoCRR:=b#N#W0H8El5LFR8,L8IHC
2;
FSOMN#0MM0RC_C8bCHbL#kVRH:RMo0CC:sR=CRMC08_FH_bbHCDMNC5I0H8EL,RI0H8E
2;
HS#oDMNRRC4RRRRR#:R0D8_FOoH_OPC05Fs4FR8IFM0R;j2
HS#oDMNRRC.RRRRR#:R0D8_FOoH_OPC05Fs4FR8IFM0R;j2
SSSSRSR
RRR#MHoNqDR0lsHR:RRR8#0_oDFHPO_CFO0sI5NH-8C4FR8IFM0R;j2
RRR#MHoNADR0lsHR:RRR8#0_oDFHPO_CFO0sI5LH-8C4FR8IFM0R;j2
R
RRo#HMRNDqHbslRCR:0R#8F_Do_HOP0COFNs5I-H84FR8IFM0R;j2
RRR#MHoNADRblsHC:RRR8#0_oDFHPO_CFO0sI5LH48-RI8FMR0Fj
2;R#RRHNoMDER1Fus0RRR:#_08DHFoOC_POs0F5HNI8I+LH48-RI8FMR0Fj:2R=FR50sEC#>R=R''j2
;
R#RRHNoMDCR)#0kD4RR:#_08DHFoOC_POs0F5HNI8LC+ICH8-84RF0IMF2Rj;R
RRo#HMRND)kC#DR0G:0R#8F_Do_HOP0COFNs5ICH8+HLI84C-RI8FMR0Fj
2;R#RRHNoMDCR)#0kDNRR:#_08DHFoOC_POs0F5HNI8LC+ICH8-84RF0IMF2Rj;R
RRo#HMRND)kC#DR0L:0R#8F_Do_HOP0COFNs5ICH8+HLI84C-RI8FMR0Fj
2;R#RRHNoMDCR)#0kDCRR:#_08DHFoOC_POs0F5HNI8LC+ICH8-84RF0IMF2Rj;R

RHR#oDMNRFus8R4,u8sF4k_NGu,Rs4F8_#sCR:RRR8#0_oDFHPO_CFO0sI5NH+8CL8IHCR-48MFI0jFR2R;
RHR#oDMNRFus8R.RR#:R0D8_FOoH_OPC05FsI0H8ER-48MFI0jFR2
;
SlOFbCFMMe0R.mApBSi
SMoCCOsHRS5
SISNHE80RH:RMo0CC:sR=IRNH
8;SLSSI0H8ERR:HCM0oRCs:L=RI;H8
SSSM8CC_bbHCVLk#RR:HCM0o2Cs;S
Sb0FsRS5
SRSqR:RRRRHMR8#0_oDFHPO_CFO0sI5NH48-RI8FMR0Fj
2;SASSRRRR:MRHR0R#8F_Do_HOP0COFLs5I-H84FR8IFM0R;j2
SSSu7)mRF:Rk#0R0D8_FOoH_OPC05FsN8IH+HLI8R-48MFI0jFR2
2;S8CMRlOFbCFMM
0;
oLCHRMR-L-RD	FO_Dlk0S

-b-RkFsb#RC:0CN	RsONCVRFRC0ERN4RM.8R-0LHR#ONCS#
-0-R$RbCRRR:OLFlH0MNHNFMD-
S-MRHb#k0Rq:R,
RASR--Fbk0k:0#Rmu)7-
S-sR0H0lREHCRM0bk#FR0RRLCMIFRHs8CRN0EMER0CkRF00bk
VSH_bbHCR4:H5VRM8CC_bbHCVLk#RR=4o2RCsMCN
0CSsS0H0lH_Rq:VRFsHMRHR0jRFIRNH-8C4CRoMNCs0SC
S0SN0LsHkR0C\N3sMR	\FsVRCqo#RD:RNDLCRRH#jS;
S0SN0LsHkR0C\F3b8\ClRRFVs#CoqRR:DCNLD#RHR
H;SNSS0H0sLCk0Rb\3Fl8CL\k#RRFVs#CoqRR:DCNLD#RHR""q;S
SS0N0skHL0\CR38lFk\DCRRFVs#CoqRR:DCNLD#RHRv"1z"pa;S
SS0N0skHL0\CR3lsCF_PCMIF_N\sMRRFVs#CoqRR:DCNLD#RHR
4;SCSLo
HMSsSSCqo#:bRRHLbCkSV
SFSbsl0RN
b5SSSSS=QR>5RqH
2,SSSSS=mR>0Rqs5HlH;22
CSSMo8RCsMCNR0C0lsHHq0_;S

SH0slAH0:FRVsRRHHjMRRR0FL8IHCR-4oCCMsCN0
SSSNs00H0LkC3R\s	NM\VRFRosC#:ARRLDNCHDR#;Rj
SSSNs00H0LkC3R\bCF8lF\RVCRsoR#A:NRDLRCDHH#R;S
SS0N0skHL0\CR38bFCklL#F\RVCRsoR#A:NRDLRCDH"#RA
";SNSS0H0sLCk0Rl\3FD8kCF\RVCRsoR#A:NRDLRCDH"#R1pvza
";SNSS0H0sLCk0Rs\3CPlFCF_M_sINMF\RVCRsoR#A:NRDLRCDH4#R;S
SLHCoMS
SSosC#RA:RbbHCVLk
SSSSsbF0NRlbS5
SSSSS=QR>5RAH
2,SSSSSRSm=A>R0lsH52H2;S
SCRM8oCCMsCN0RH0slAH0;C
SMo8RCsMCNR0CHbV_H4bC;H
SVH_bb:CjRRHV5CMC8H_bbkCLV=#RRRj2oCCMsCN0
qSS0lsHRR<=qI5NH-8C4FR8IFM0R;j2
ASS0lsHRR<=AI5LH-8C4FR8IFM0R;j2
MSC8CRoMNCs0HCRVH_bb;Cj
-
S-CRslCFPRC0ER0CGsLNRHR0#N00REpCR1CARMR8
RsRbkHMC0b:RsCFO#5#RqH0slA,R0lsH2L
SCMoHR-R-RFbsO#C#RkbsM0CH
HSSVlRNF=8RR04RE
CMSCSS4=R<R''jRq&R0lsH5;j2
SSSqHbsl<CR=0Rqs5HlN8IHCR-48MFI04FR2S;
S#CDHNVRlRF8=RR.0MEC
RRRRRRRR4RCRR<=qH0slR548MFI0jFR2S;
SbSqsCHlRR<=qH0slI5NH-8C4FR8IFM0R;.2
RRRRCRRD
#CSCSS4=R<R''jR'&Rj
';SqSSblsHC=R<Rsq0H
l;SMSC8VRH;S

SRHVL8lFR4=RRC0EMS
SSRC.<'=Rj&'RRsA0Hjl52S;
SbSAsCHlRR<=AH0slI5LH-8C4FR8IFM0R;42
CSSDV#HRFLl8RR=.ER0CRM
RRRRRRRRC<.R=0RAs5Hl4FR8IFM0R;j2
SSSAHbsl<CR=0RAs5HlL8IHCR-48MFI0.FR2R;
RRRRR#CDCS
SSRC.<'=Rj&'RR''j;S
SSsAbHRlC<A=R0lsH;S
SCRM8H
V;S8CMRFbsO#C#RkbsM0CH;S

-v-RkHD0bRD$L0$RECCRGN0sR0LH#VRHRRICECNPRCFMRRFs0RIFCsG0NHRL0F#RV
RqS_HVNR4:H5VRN8lF=R42oCCMsCN0
HSSV4_NLRj:H5VRL8lFRR<=jsRFRFLl8RR>.o2RCsMCN
0CS)SSCD#k0<NR=mRBh1e_ap7_mBtQ_Be a5m)jN,RICH8+HLI8RC2IMECR45C5Rj2=jR''
2RSSSSSRSRCCD#Ra1X5sAbH,lCRHNI8LC+ICH82R;
RRRRR8CMRMoCC0sNCVRH_LN4jS;
S_HVN44L:VRHRl5LF=8RRR42oCCMsCN0
SSS)kC#DR0N<B=Rm_he1_a7pQmtB _eB)am5Rj,N8IHCI+LH28CRCIEMCR5425jR'=RjR'2
SSSSRSSR#CDCXR1ab5AsCHlR'&RjR',N8IHCI+LH28C;R
RRRRRCRM8oCCMsCN0R_HVN44L;S
SHNV_4:L.RRHV5FLl8RR=.o2RCsMCN
0CS)SSCD#k0<NR=mRBh1e_ap7_mBtQ_Be a5m)jN,RICH8+HLI8RC2IMECR45C5Rj2=jR''
2RSSSSSRSRCCD#Ra1X5sAbHRlC&jR''RR&',j'RHNI8LC+ICH82R;
RRRRR8CMRMoCC0sNCVRH_LN4.S;
CRM8oCCMsCN0R_HVN
4;SNHVMR.:H5VRN8lF=N.RMN8RI0H8E2>.RMoCC0sNC-RR-hRz1hQt R7
RRRRRo#HMRNDMEF1H,V0RH#EV80C,8RN8RC8:0R#8F_Do_HOP0COFNs5ICH8+HLI84C-RI8FMR0Fj
2;SoLCHSM
SNHVMj.L:VRHRl5LF<8R=RRjFLsRlRF8>2R.RMoCC0sNCR
RRMSSFH1EV<0R=XR1ab5AsCHl,IRNH+8CL8IHC
2;RRRRRMRC8CRoMNCs0HCRV.NML
j;SVSHNLM.4H:RVLR5lRF8=2R4RMoCC0sNCR
RRMSSFH1EV<0R=XR1ab5AsCHlR'&RjR',N8IHCI+LH28C;R
RRRRRCRM8oCCMsCN0RNHVM4.L;S
SHMVN.:L.RRHV5FLl8RR=.o2RCsMCN
0CRSRRS1MFE0HVRR<=15XaAHbsl&CRR''jR'&RjR',N8IHCI+LH28C;R
RRRRRCRM8oCCMsCN0RNHVM..L;S
S#VEH0RC8<M=RFH1EVN05ICH8+HLI8.C-RI8FMR0Fj&2RR''j;R
RRRRRNC888RRR<M=RFH1EV+0RRH#EV80C;S
S)kC#DR0N<B=Rm_he1_a7pQmtB _eB)am5Nj,ICH8+HLI8RC2IMECR45CR"=Rj2j"
SSSSRSRCCD#R1MFE0HVRCIEMCR54RR=""j42S
SSRSSR#CDCER#HCV08ERIC5MRC=4RRj"4"S2
SSSSRDRC#NCR888C;-SR-5RRC=4RR4"4"S2
CRM8oCCMsCN0RNHVM
.;S_HVNR.:H5VRN8lF=N.RMN8RI0H8E2=.RMoCC0sNC-RR-QR1t7h 
#SSHNoMDFRM1VEH0O,RFDlbCMlC00,RIFFOl:bRR8#0_oDFHPO_CFO0sI5NH+8CL8IHCR-48MFI0jFR2S;
LHCoMS
SHNV_.:LjRRHV5FLl8=R<RFjRslRLF>8RRR.2oCCMsCN0
RRRRMSSFH1EV<0R=XR1ab5AsCHl,IRNH+8CL8IHC
2;RRRRRMRC8CRoMNCs0HCRV._NL
j;SVSH_LN.4H:RVLR5lRF8=2R4RMoCC0sNCR
RRMSSFH1EV<0R=XR1ab5AsCHlR'&RjR',N8IHCI+LH28C;R
RRRRRCRM8oCCMsCN0R_HVN4.L;S
SHNV_.:L.RRHV5FLl8RR=.o2RCsMCN
0CRSRRS1MFE0HVRR<=15XaAHbsl&CRR''jR'&RjR',N8IHCI+LH28C;R
RRRRRCRM8oCCMsCN0R_HVN..L;S
SObFlDCClM<0R=FRM0FRM1VEH0S;
SF0IObFlRR<=ObFlDCClM+0RR''4;R
RRRRR)kC#DR0N<B=Rm_he1_a7pQmtB _eB)am5Rj,N8IHCI+LH28CRCIEMCR54RR=""jj2S
SSRSSR#CDCFRM1VEH0ERIC5MRC=4RR4"j"S2
SSSSRDRC#0CRIFFOlIbRERCM5RC4=4R"4
"2SSSSSCRRDR#C0OIFF5lbN8IHCI+LH-8C.FR8IFM0RRj2&jR''R;R-I-RERCM5RC4=4R"j
"2S8CMRMoCC0sNCVRH_;N.
-
S-kRvDb0HDL$R$ER0CGRC0RsNL#H0RRHVIECRNRPCFRMCF0sRICFRGN0sR0LH#VRFRSA
HLV_4H:RVLR5l=F84o2RCsMCN
0CRRRRRVRH_NL4jR:RH5VRN8lFRR<=jsRFRFNl8RR>.o2RCsMCN
0CS)SSCD#k0<LR=mRBh1e_ap7_mBtQ_Be a5m)jN,RICH8+HLI8RC2IMECR.5C5Rj2=jR''
2RSSSSSRSRCCD#Ra1X5sqbH,lCRHNI8LC+ICH82R;
RRRRR8CMRMoCC0sNCVRH_NL4jS;
S_HVL44N:VRHRl5NF=8RRR42oCCMsCN0
SSS)kC#DR0L<B=Rm_he1_a7pQmtB _eB)am5Rj,N8IHCI+LH28CRCIEMCR5.25jR'=RjR'2
SSSSRSSR#CDCXR1ab5qsCHlR'&RjR',N8IHCI+LH28C;R
RRRRRCRM8oCCMsCN0R_HVL44N;S
SHLV_4:N.RRHV5FNl8RR=.o2RCsMCN
0CS)SSCD#k0<LR=mRBh1e_ap7_mBtQ_Be a5m)jN,RICH8+HLI8RC2IMECR.5C5Rj2=jR''
2RSSSSSRSRCCD#Ra1X5sqbHRlC&jR''RR&',j'RHNI8LC+ICH82R;
RRRRR8CMRMoCC0sNCVRH_NL4.S;
CRM8oCCMsCN0R_HVL
4;RHRRV.LM:VRHRl5LF.8=R8NMRHLI8>0E.o2RCsMCNR0CRR--zQh1t7h 
RRRR#RRHNoMDFRM1VEH0#,RE0HVCR8,NC888RR:#_08DHFoOC_POs0F5HNI8LC+ICH8-84RF0IMF2Rj;L
SCMoH
HSSV.LMNRj:H5VRN8lFRR<=jsRFRFNl8RR>.o2RCsMCN
0CRSRRS1MFE0HVRR<=15XaqHbslRC,N8IHCI+LH28C;R
RRRRRCRM8oCCMsCN0RLHVMj.N;S
SHMVL.:N4RRHV5FNl8RR=4o2RCsMCN
0CRSRRS1MFE0HVRR<=15XaqHbsl&CRR''j,IRNH+8CL8IHC
2;RRRRRMRC8CRoMNCs0HCRV.LMN
4;SVSHLNM..H:RVNR5lRF8=2R.RMoCC0sNCR
RRMSSFH1EV<0R=XR1ab5qsCHlR'&Rj&'RR''j,IRNH+8CL8IHC
2;RRRRRMRC8CRoMNCs0HCRV.LMN
.;SES#HCV08=R<R1MFE0HV5HNI8LC+ICH8-8.RF0IMF2RjR'&Rj
';RRRRR8RN8RC8R=R<R1MFE0HVR#+RE0HVC
8;SCS)#0kDL=R<RhBmea_17m_pt_QBea Bmj)5,IRNH+8CL8IHCI2RERCM5RC.=jR"j
"2SSSSSCRRDR#CMEF1HRV0IMECR.5CR"=Rj24"
SSSSRSRCCD#RH#EV80CRCIEMCR5.RR=""4j2S
SSRSSR#CDC8RN8;C8R-RR-5RRC=.RR4"4"S2
CRM8oCCMsCN0RLHVM
.;S_HVLR.:H5VRL8lF=N.RML8RI0H8E2=.RMoCC0sNC-RR-QR1t7h 
#SSHNoMDFRM1VEH0O,RFDlbCMlC00,RIFFOl:bRR8#0_oDFHPO_CFO0sI5NH+8CL8IHCR-48MFI0jFR2S;
LHCoMR
RRRRRHLV_.:NjRVRHRl5NF<8R=RRjFNsRlRF8>2R.RMoCC0sNCR
RRRRRRMRRFH1EV<0R=XR1ab5qsCHl,IRNH+8CL8IHC
2;SMSC8CRoMNCs0HCRV._LN
j;SVSH_NL.4H:RVNR5lRF8=2R4RMoCC0sNCR
RRMSSFH1EV<0R=XR1ab5qsCHlR'&RjR',N8IHCI+LH28C;R
RRRRRCRM8oCCMsCN0R_HVL4.N;S
SHLV_.:N.RRHV5FNl8RR=.o2RCsMCN
0CRSRRS1MFE0HVRR<=15XaqHbsl&CRR''jR'&RjR',N8IHCI+LH28C;R
RRRRRCRM8oCCMsCN0R_HVL..N;S
SObFlDCClM<0R=FRM0FRM1VEH0S;
SF0IObFlRR<=ObFlDCClM+0RR''4;S
S)kC#DR0L<B=Rm_he1_a7pQmtB _eB)am5Rj,N8IHCI+LH28CRCIEMCR5.RR=""jj2S
SSRSSR#CDCFRM1VEH0ERIC5MRC=.RR4"j"S2
SSSSRDRC#0CRIFFOlIbRERCM5RC.=4R"4
"2SSSSSCRRDR#C0OIFF5lbN8IHCI+LH-8C4FR8IFM0RRj2&jR''R;R-I-RERCM5RC.=4R"j
"2S8CMRMoCC0sNCVRH_;L.
-
S-kRvDb0HD0$RECCRGN0sR0LH#VRHRRICECNPR0CGsRN#HCMRHC0EsRRqNRM8AH
SV#_C:VRHRN55lRF8=RR4FNsRlRF8=2R.R8NMRl5LF=8RRF4RslRLF=8RR2.2RMoCC0sNCS
S)kC#D50Cd<2R=CRR4254R8NMR5C4jN2RMC8R.254R8NMR5C.j
2;SCS)#0kDC25.RR<=55C44N2RM58RMRF0Cj452N2RMC8R.2542sRF
SSSSRSSR45C5R42NRM8C4.52MRN8MR5FC0R.25j2
2;SCS)#0kDC254RR<=55C44N2RM58RMRF0Cj452N2RMC8R.25j2sRF
SSSSRSSRM55FC0R42542MRN84RC5Rj2NRM8C4.52F2RsS
SSSSSRCR54254R8NMRF5M0.RC5242R8NMR5C.jR22FSs
SSSSS5RRCj452MRN8.RC5R42NRM850MFR5C.j222;S
S)kC#D50Cj<2R=CRR425jR8NMR5C.j
2;SVSH_#sCCH:RVNR5ICH8+HLI8>CRRRc2oCCMsCN0
SSS)kC#D50CN8IHCI+LH-8C4FR8IFM0RRc2<B=Rm_he1_a7pQmtB _eB)am5Rj,N8IHCI+LHR8C-2Rc;S
SCRM8oCCMsCN0R_HVsCC#;C
SMo8RCsMCNR0CHCV_#
;
SkLlDR0:HNVRICH8R.>RR8NMRHLI8>CRRo.RCsMCN
0CSkSlDG0GRe:R.mApBSi
SCSoMHCsONRlb
R5SSSSSISNHE80RR=>N8IH,S
SSSSSL8IH0=ER>IRLH
8,SSSSSCSMCb8_HLbCkRV#=M>RC_C8bCHbL#kV2S
SSsbF0NRlb
R5SSSSSRqRR>R=RsqbH,lC
SSSSRSAR=RR>bRAsCHl,S
SSuSS)Rm7=1>RE0Fsu
2;S8CMRMoCC0sNClRLk;D0
R
RR0CGCHM80b:RsCFO#5#R1sEF0
u2SoLCHRMR-b-RsCFO#C#RGM0C8
H0RRRRRCR)#0kD4=R<Ra1X5F1Es,0uRHNI8LC+ICH82S;
CRM8bOsFCR##CCG0M08H;R

RLRNljF8:VRHRN55l>F8.sRFRFNl82=jR8NMRl5LF.8>RRFsL8lF=2j2RMoCC0sNCS
S)kC#DR0G<)=RCD#k0
4;S8CMRMoCC0sNCLRNljF8;R

RLRNl4F8:VRHRl5NF48=R8NMRl5LF.8>RRFsL8lF=2j2RRFs5l5NF.8>RRFsN8lF=Rj2NRM8L8lF=R42oCCMsCN0
)SSCD#k0<GR=CR)#0kD4I5NH+8CL8IHCR-.8MFI0jFR2RR&';j'
MSC8CRoMNCs0NCRL8lF4
;
RNRRL8lF.H:RVNR5l=F84MRN8lRLF48=2sRFRl5NF.8=R8NMRl5LF.8>RRFsL8lF=2j2RRFs5l5NF.8>RRFsN8lF=Rj2NRM8L8lF=R.2oCCMsCN0
)SSCD#k0<GR=CR)#0kD4I5NH+8CL8IHCR-d8MFI0jFR2RR&""jj;C
SMo8RCsMCNR0CNFLl8
.;
RRRNFLl8Rd:H5VRN8lF=N.RML8Rl=F84F2RsNR5l=F84MRN8lRLF.8=2CRoMNCs0SC
S#)CkGD0RR<=)kC#D504N8IHCI+LH-8CcFR8IFM0RRj2&jR"j;j"
MSC8CRoMNCs0NCRL8lFd
;
RNRRL8lFcH:RVNR5l=F8.MRN8lRLF.8=2CRoMNCs0SC
S#)CkGD0RR<=)kC#D504N8IHCI+LH-8C6FR8IFM0RRj2&jR"j"jj;C
SMo8RCsMCNR0CNFLl8
c;
HRSVC_oMNCs0RC:H5VR5l5NF>8RRRj2NRM85FNl8RR<dR22F5sR5FLl8RR>jN2RM58RL8lFRd<R2R22oCCMsCN0
RRRLHCoMS
SH#V_0CN04H:RV5R5N8lFRj>R2MRN8NR5lRF8<2RdR8NMRl5LF>8RRRj2NRM85FLl8RR<dR22oCCMsCN0
SSSu8sF4k_NG=R<RCR)#0kDNRR+)kC#DR0L+CR)#0kDCS;
S8CMRMoCC0sNCVRH_N#00;C4
HSSV0_#N.0C:VRHRN55lRF8>2RjR8NMRl5NF<8RRRd2NRM85l5LF>8RRR.2F5sRL8lFRj=R2R22oCCMsCN0
SSSu8sF4k_NG=R<RCR)#0kDNS;
S8CMRMoCC0sNCVRH_N#00;C.
HSSV0_#Nd0C:VRHRL55lRF8>2RjR8NMRl5LF<8RRRd2NRM85l5NF>8RRR.2F5sRN8lFRj=R2R22oCCMsCN0
SSSu8sF4k_NG=R<RCR)#0kDLS;
S8CMRMoCC0sNCVRH_N#00;Cd
S
SHbV_H4bN:VRHRC5MCb8_HLbCkRV#=2R4RMoCC0sNCS
SSbbHCRj:VRFsHMRHR0jRFHRI8-0E4CRoMNCs0SC
SNSS0H0sLCk0Rs\3N\M	RRFVs#Co1RR:DCNLD#RHR
4;SSSSNs00H0LkC3R\LHCoMs_0CRC\FsVRC1o#RD:RNDLCRRH#4S;
SNSS0H0sLCk0Rs\3CPlFCF_M_sINMF\RVCRsoR#1:NRDLRCDH4#R;S
SSoLCHSM
SsSSC1o#:bRRHLbCkSV
SbSSFRs0l5Nb
SSSSQSSRR=>u8sF4k_NG25H,S
SSSSSm>R=RFus8s4_CH#52
2;SCSSMo8RCsMCNR0CbCHbjS;
S8CMRMoCC0sNCVRH_bbHN
4;SVSH_bbHNRj:H5VRM8CC_bbHCVLk#RR=jo2RCsMCN
0CSuSSs4F8_#sCRR<=u8sF4k_NGS;
S8CMRMoCC0sNCVRH_bbHN
j;S8CMRMoCC0sNCVRH_MoCC0sNC
;
RVSH_MoCC0sNC:_4RRHV5l5NF>8RRR.2NRM85FLl8RR>.R22oCCMsCN0
uSSs4F8_#sCRR<=RhBmea_17m_pt_QBea Bmj)5,IRNH+8CL8IHC
2;S8CMRMoCC0sNCVRH_MoCC0sNC;_4
R
RRFus8<4R=CR)#0kDGRR+u8sF4C_s#
;
S0CGCbM8s:F8RFbsO#C#Rs5uF284
CSLoRHMRR--bOsFCR##CCG0Ms8bFS8
SRHVI0H8ERR>N8IHCRR+L8IHCER0CSM
SsSuFR8.<1=RXua5s4F8,HRI820E;S
SCCD#
SSSu8sF.=R<RFus8I45HE80-84RF0IMF2Rj;S
SCRM8H
V;S8CMRFbsO#C#R0CGCbM8s;F8
H
SVH_bb:L4RRHV5CMC8H_bbkCLV=#RRR42oCCMsCN0
LSSkkVF00bk:FRVsRRHHjMRRR0FI0H8ER-4oCCMsCN0
SSSNs00H0LkC3R\s	NM\VRFRosC#:1RRLDNCHDR#;R.
SSSNs00H0LkC3R\C_M80CsC\VRFRosC#:1RRLDNCHDR#;R4
SSSNs00H0LkC3R\bCF8lF\RVCRsoR#1:NRDLRCDHH#R;S
SS0N0skHL0\CR38bFCklL#F\RVCRsoR#1:NRDLRCDH"#Ru7)m"S;
S0SN0LsHkR0C\C3slCFP__MFIMNs\VRFRosC#:1RRLDNCHDR#;R4
LSSCMoH
SSSs#Co1R:RbCHbL
kVSSSSSsbF0NRlbS5
SSSSSRSQ=u>Rs.F85,H2
SSSSSSSm>R=Rmu)725H2S;
S8CMRMoCC0sNCkRLV0Fkb;k0
MSC8CRoMNCs0HCRVH_bb;L4
VSH_bbHLRj:H5VRM8CC_bbHCVLk#RR=jo2RCsMCN
0CS)Sum<7R=sRuF;8.
MSC8CRoMNCs0HCRVH_bb;Lj
M
C8DRLF_O	l0kD;



