library verilog;
use verilog.vl_types.all;
entity dffprqnx4v1mce is
    port(
        CDN             : in     vl_logic;
        CK              : in     vl_logic;
        D               : in     vl_logic;
        Q               : out    vl_logic;
        QN              : out    vl_logic
    );
end dffprqnx4v1mce;
