library verilog;
use verilog.vl_types.all;
entity dp_spare_gate is
    port(
        signal_in       : in     vl_logic
    );
end dp_spare_gate;
