library verilog;
use verilog.vl_types.all;
entity cfg_cntl is
    port(
        ctrl_sfdp_en    : out    vl_logic;
        njbse_sign_read : out    vl_logic;
        njbse_sign_cmd  : out    vl_logic;
        njbse_sign_cmd_read: out    vl_logic;
        ctrl_smfreq_sel : out    vl_logic_vector(1 downto 0);
        jtag_active_smsync: out    vl_logic;
        jtag_active_smsync_jb: out    vl_logic;
        buf128_dat      : out    vl_logic_vector(127 downto 0);
        sector_dat      : out    vl_logic_vector(15 downto 0);
        sector_erase    : out    vl_logic_vector(11 downto 0);
        ctrl0           : out    vl_logic_vector(31 downto 0);
        ctrl1           : out    vl_logic_vector(31 downto 0);
        sd_trim         : out    vl_logic_vector(255 downto 0);
        cfg_i2c_dat     : out    vl_logic_vector(15 downto 0);
        isc_exec_a      : out    vl_logic;
        isc_exec_b      : out    vl_logic;
        isc_exec_c      : out    vl_logic;
        isc_exec_d      : out    vl_logic;
        isc_exec_e      : out    vl_logic;
        isc_exec_f      : out    vl_logic;
        fl_erase_exec   : out    vl_logic;
        gsrn            : out    vl_logic;
        gsrn_sync       : out    vl_logic;
        goe             : out    vl_logic;
        ts_all          : out    vl_logic;
        done_gwe        : out    vl_logic;
        freeze_io       : out    vl_logic;
        freeze_mib      : out    vl_logic;
        pcs_rstn        : out    vl_logic;
        en_pupn         : out    vl_logic;
        isc_operational : out    vl_logic;
        isc_disable_exec: out    vl_logic;
        sed_rst_async   : out    vl_logic;
        sed_rst_sync    : out    vl_logic;
        sed_rst_flag    : out    vl_logic;
        cfg_sed_en      : out    vl_logic;
        dev_sed_exec    : out    vl_logic;
        fl_start_ppt    : out    vl_logic;
        fl_start_cdm    : out    vl_logic;
        fl_start_sdm0   : out    vl_logic;
        fl_start_sdm1   : out    vl_logic;
        fl_start_sdm2   : out    vl_logic;
        fl_start_sdm_cfg0: out    vl_logic;
        fl_start_sdm_cfg1: out    vl_logic;
        authdone_sdm0_start: out    vl_logic;
        authdone_sdm1_start: out    vl_logic;
        access_flash_all: out    vl_logic;
        access_sudo     : out    vl_logic;
        start_bke       : out    vl_logic;
        ebr_init_en     : out    vl_logic;
        dev_sdm_cfg0_exec: out    vl_logic;
        dev_sdm_cfg1_exec: out    vl_logic;
        finish_bse      : out    vl_logic;
        fail_bse        : out    vl_logic;
        busy_bse        : out    vl_logic;
        comp_dic        : out    vl_logic_vector(127 downto 0);
        initn_tmr       : out    vl_logic;
        goe_tmr         : out    vl_logic;
        done_tmr        : out    vl_logic;
        ref_boot0       : out    vl_logic;
        ref_boot1       : out    vl_logic;
        ref_boot2       : out    vl_logic;
        isc_rst_async   : out    vl_logic;
        isc_rst_sync    : out    vl_logic;
        sf_rst_async    : out    vl_logic;
        sf_rst_sync     : out    vl_logic;
        nj_rst_async    : out    vl_logic;
        nj_rst_sync0    : out    vl_logic;
        nj_rst_sync     : out    vl_logic;
        nji2c_rst_async : out    vl_logic;
        njtrx_rst_async : out    vl_logic;
        njtrx_rst_async0: out    vl_logic;
        restart_bse_en  : out    vl_logic;
        njboot_dat      : out    vl_logic_vector(7 downto 0);
        cfg_mstr_start  : out    vl_logic;
        cfg_mstr_stop   : out    vl_logic;
        cfg_mtx_dat     : out    vl_logic_vector(7 downto 0);
        cfg_mcsn_dat    : out    vl_logic_vector(7 downto 0);
        ref_launch      : out    vl_logic;
        ref_sys_slow    : out    vl_logic;
        njbse_preamble  : out    vl_logic;
        njbse_sstcmd    : out    vl_logic;
        njbse_txcmd     : out    vl_logic;
        njbse_rxcmd     : out    vl_logic;
        njbse_rxdec     : out    vl_logic;
        njbse_rxall     : out    vl_logic;
        njbse_bypass    : out    vl_logic;
        njbse_fthrough  : out    vl_logic;
        tx_setmcpu      : out    vl_logic;
        tx_command      : out    vl_logic;
        tx_operand      : out    vl_logic;
        fsd_persistn_progn: out    vl_logic;
        fsd_persist_initn: out    vl_logic;
        fsd_persist_done: out    vl_logic;
        fsd_persistn_jtag: out    vl_logic;
        fsd_persistn_sspi: out    vl_logic;
        fsd_persistn_i2c: out    vl_logic;
        fsd_persist_mspi: out    vl_logic;
        fsd_boot_sel    : out    vl_logic_vector(2 downto 0);
        sd_i2c_addr     : out    vl_logic_vector(7 downto 0);
        cib_wkupclk_en  : out    vl_logic;
        cfg_ctrl0_upd   : out    vl_logic;
        j_com_word4_dat : out    vl_logic_vector(127 downto 0);
        nj_com_word4_dat: out    vl_logic_vector(127 downto 0);
        jinstr_cap      : out    vl_logic_vector(7 downto 0);
        jconfig_cap     : out    vl_logic_vector(7 downto 0);
        jburst_inp      : out    vl_logic;
        dryrun_inp      : out    vl_logic;
        busy_int        : out    vl_logic;
        ref_exit        : out    vl_logic;
        instr_dts       : out    vl_logic;
        start_dts       : out    vl_logic;
        last_addr_cib   : out    vl_logic_vector(15 downto 0);
        cfg_done_cib    : out    vl_logic;
        busy_seldr      : out    vl_logic;
        isc_done        : out    vl_logic;
        lsc_done        : out    vl_logic;
        lsc_done_ebr    : out    vl_logic;
        lsc_done_ip     : out    vl_logic;
        lsc_done_hse    : out    vl_logic;
        wkup_done       : out    vl_logic;
        mfg_margin_en   : out    vl_logic;
        exit_accessed   : out    vl_logic;
        isc_data_shift_iqual: out    vl_logic;
        lsc_prog_incr_rti_iqual: out    vl_logic;
        lsc_prog_incr_enc_iqual: out    vl_logic;
        lsc_prog_incr_cmp_iqual: out    vl_logic;
        lsc_prog_incr_cne_iqual: out    vl_logic;
        isc_data_shift_cqual: out    vl_logic;
        lsc_prog_incr_rti_cqual: out    vl_logic;
        lsc_prog_incr_enc_cqual: out    vl_logic;
        lsc_prog_incr_cmp_cqual: out    vl_logic;
        lsc_prog_incr_cne_cqual: out    vl_logic;
        cfg_reset_crc16 : out    vl_logic;
        lsc_reboot_cq   : out    vl_logic;
        lsc_read_pes_qual: out    vl_logic;
        sf_prog_ucode_qual: out    vl_logic;
        sf_program_qual : out    vl_logic;
        sf_read_qual    : out    vl_logic;
        sf_erase_qual   : out    vl_logic;
        sf_prog_done_qual: out    vl_logic;
        sf_erase_done_qual: out    vl_logic;
        sf_prog_sec_qual: out    vl_logic;
        sf_init_addr_qual: out    vl_logic;
        sf_write_addr_qual: out    vl_logic;
        sf_address_shift_qual: out    vl_logic;
        sf_prog_incr_rti_qual: out    vl_logic;
        sf_prog_incr_enc_qual: out    vl_logic;
        sf_prog_incr_cmp_qual: out    vl_logic;
        sf_prog_incr_cne_qual: out    vl_logic;
        sf_vfy_incr_rti_qual: out    vl_logic;
        sf_prog_sed_crc_qual: out    vl_logic;
        sf_read_sed_crc_qual: out    vl_logic;
        sf_write_bus_addr_qual: out    vl_logic;
        sf_pcs_write_qual: out    vl_logic;
        sf_pcs_read_qual: out    vl_logic;
        sf_ebr_write_qual: out    vl_logic;
        sf_ebr_read_qual: out    vl_logic;
        sf_prog_sec_eqv : out    vl_logic;
        sed_init_addr_qual: out    vl_logic;
        sed_write_addr_qual: out    vl_logic;
        sed_read_incr_qual: out    vl_logic;
        sed_prog_sed_crc_qual: out    vl_logic;
        fl_prog_ucode_qual: out    vl_logic;
        fl_prog_done_qual: out    vl_logic;
        fl_prog_sec_qual: out    vl_logic;
        fl_prog_secplus_qual: out    vl_logic;
        fl_disable_done0_qual: out    vl_logic;
        fl_disable_done1_qual: out    vl_logic;
        fl_erase_qual   : out    vl_logic;
        fl_erase_all_qual: out    vl_logic;
        fl_init_addr_qual: out    vl_logic;
        fl_write_addr_qual: out    vl_logic;
        fl_prog_incr_nv_qual: out    vl_logic;
        fl_read_incr_nv_qual: out    vl_logic;
        fl_prog_password_qual: out    vl_logic;
        fl_prog_cipher_key0_qual: out    vl_logic;
        fl_prog_cipher_key1_qual: out    vl_logic;
        fl_prog_feature_qual: out    vl_logic;
        fl_prog_feabits_qual: out    vl_logic;
        fl_init_addr_ufm_qual: out    vl_logic;
        fl_prog_tag_qual: out    vl_logic;
        fl_erase_tag_qual: out    vl_logic;
        fl_read_tag_qual: out    vl_logic;
        fl_prog_pes_qual: out    vl_logic;
        fl_prog_mes_qual: out    vl_logic;
        fl_prog_hes_qual: out    vl_logic;
        fl_prog_trim0_qual: out    vl_logic;
        fl_prog_trim1_qual: out    vl_logic;
        fl_read_hes_qual: out    vl_logic;
        fl_prog_csec_qual: out    vl_logic;
        fl_prog_usec_qual: out    vl_logic;
        fl_prog_uds_qual: out    vl_logic;
        fl_udss0_authdone_exec: out    vl_logic;
        fl_udss1_authdone_exec: out    vl_logic;
        fl_prog_authmode_qual: out    vl_logic;
        fl_prog_aesfea_qual: out    vl_logic;
        fl_mtest_qual   : out    vl_logic;
        mfg_flash_en    : out    vl_logic;
        stdby_ena       : out    vl_logic;
        dev_stdby_exec  : out    vl_logic;
        dev_sleep_exec  : out    vl_logic;
        dev_wkup_exec   : out    vl_logic;
        lsc_i2ci_crbr_wt_qual: out    vl_logic;
        lsc_i2ci_txdr_wt_qual: out    vl_logic;
        lsc_i2ci_rxdr_rd_qual: out    vl_logic;
        lsc_i2ci_sr_rd_qual: out    vl_logic;
        lsc_auth_ctrl_cqual: out    vl_logic;
        key_byte        : out    vl_logic_vector(7 downto 0);
        sd_aes_key      : out    vl_logic_vector(255 downto 0);
        sd_auth_en      : out    vl_logic_vector(1 downto 0);
        sd_rand_noise   : out    vl_logic;
        sd_rand_aes     : out    vl_logic;
        finish_cdm      : out    vl_logic;
        fl_prog_pubkey0_qual: out    vl_logic;
        fl_prog_pubkey1_qual: out    vl_logic;
        fl_prog_pubkey2_qual: out    vl_logic;
        fl_prog_pubkey3_qual: out    vl_logic;
        sd_authdone_cfg0: out    vl_logic;
        sd_authdone_cfg1: out    vl_logic;
        sd_sec_jtag     : out    vl_logic_vector(1 downto 0);
        sd_sec_sspi     : out    vl_logic_vector(1 downto 0);
        sd_sec_si2c     : out    vl_logic_vector(1 downto 0);
        sd_sec_bspi     : out    vl_logic;
        sd_sec_bi2c     : out    vl_logic;
        secJTAGByCIB    : out    vl_logic;
        secSSPIByCIB    : out    vl_logic;
        secI2CByCIB     : out    vl_logic;
        cfg0_latter     : out    vl_logic;
        mem_bist_en     : out    vl_logic;
        sdm_done_sec_read: out    vl_logic;
        njbse_rst_flag  : out    vl_logic;
        bse_sdm_cfg0    : out    vl_logic;
        bse_sdm_cfg1    : out    vl_logic;
        sd_i2c_deg      : out    vl_logic;
        sd_i2c_deg_sel  : out    vl_logic;
        lsc_bitstream_burst_qual: out    vl_logic;
        sec_read_alt_sram: out    vl_logic;
        sec_prog_alt_sram: out    vl_logic;
        cmd_altsec_sram : out    vl_logic;
        njbse_init      : out    vl_logic;
        sd_uds_trn      : out    vl_logic_vector(127 downto 0);
        uidcode         : out    vl_logic_vector(63 downto 0);
        cdm_done_por    : out    vl_logic;
        preamble_timer  : in     vl_logic_vector(3 downto 0);
        preamblePass    : in     vl_logic;
        sign_match      : in     vl_logic;
        signatureCheckEvent: in     vl_logic;
        CHIPID          : in     vl_logic_vector(7 downto 0);
        CTRL0_DEFAULT   : in     vl_logic_vector(31 downto 0);
        CTRL1_DEFAULT   : in     vl_logic_vector(31 downto 0);
        IDCODE0         : in     vl_logic_vector(31 downto 0);
        ASSP_EN         : in     vl_logic;
        HFC_EN          : in     vl_logic;
        ENC_ONLY_EN     : in     vl_logic;
        trim_idcode_msb : in     vl_logic_vector(3 downto 0);
        trim_idmsb_en   : in     vl_logic_vector(3 downto 0);
        bg_cmp_out      : in     vl_logic;
        bg_rdy          : in     vl_logic;
        proc_ring_osc   : in     vl_logic;
        dts_out         : in     vl_logic_vector(31 downto 0);
        por             : in     vl_logic;
        por_sec         : in     vl_logic;
        por_trim        : in     vl_logic;
        tck             : in     vl_logic;
        smclk           : in     vl_logic;
        smclk_scan_off  : in     vl_logic;
        hse_clk         : in     vl_logic;
        wkupclk         : in     vl_logic;
        fsafe           : in     vl_logic;
        scanen          : in     vl_logic;
        gsrn_pin_sync   : in     vl_logic;
        hfc_select_pin  : in     vl_logic;
        cfg_mstr_busy   : in     vl_logic;
        njm_tr_next     : in     vl_logic;
        njm_tr_done     : in     vl_logic;
        njm_mcpu_done   : in     vl_logic;
        preamble_std    : in     vl_logic;
        preamble_enc    : in     vl_logic;
        preamble_std_ext: in     vl_logic;
        preamble_enc_ext: in     vl_logic;
        programn_tog    : in     vl_logic;
        programn_pin_sync: in     vl_logic;
        initn_pin_sync  : in     vl_logic;
        done_pin_sync   : in     vl_logic;
        boot_setup      : in     vl_logic_vector(5 downto 0);
        cfg_i2c_dout    : in     vl_logic_vector(7 downto 0);
        wbc_active      : in     vl_logic;
        p_eboot0p       : in     vl_logic;
        p_eboot1p       : in     vl_logic;
        p_eboot1s       : in     vl_logic;
        p_eboot2p       : in     vl_logic;
        p_eboot2s       : in     vl_logic;
        p_nboot         : in     vl_logic;
        p_iboot0p       : in     vl_logic;
        p_iboot1p       : in     vl_logic;
        p_iboot1s       : in     vl_logic;
        p_iboot2p       : in     vl_logic;
        p_iboot2s       : in     vl_logic;
        p_slave         : in     vl_logic;
        p_mspi0         : in     vl_logic;
        p_mspim         : in     vl_logic;
        p_mp8           : in     vl_logic;
        p_mp16          : in     vl_logic;
        p_mspi_slow     : in     vl_logic;
        p_mspi_fast     : in     vl_logic;
        p_mspi_dual     : in     vl_logic;
        p_mspi_quad     : in     vl_logic;
        p_mp8_quad      : in     vl_logic;
        p_mp16_quad     : in     vl_logic;
        p_mspi_all      : in     vl_logic;
        p_sst           : in     vl_logic;
        p_end_bpft      : in     vl_logic;
        done_rise1      : in     vl_logic;
        cfg_crc         : in     vl_logic_vector(15 downto 0);
        njm_crc_err     : in     vl_logic;
        sed_en_adv      : in     vl_logic;
        sed_busy        : in     vl_logic;
        sed_active      : in     vl_logic;
        sed_err         : in     vl_logic;
        sed_start_bse   : in     vl_logic;
        sed_boot        : in     vl_logic;
        current_sector  : in     vl_logic_vector(11 downto 0);
        fl_load_trim0   : in     vl_logic;
        fl_load_trim1   : in     vl_logic;
        fl_load_pes     : in     vl_logic;
        fl_load_mes     : in     vl_logic;
        fl_load_pwd     : in     vl_logic;
        fl_load_fea     : in     vl_logic;
        fl_load_feabits : in     vl_logic;
        fl_load_udss0   : in     vl_logic;
        fl_load_ufs0    : in     vl_logic;
        fl_load_tss     : in     vl_logic;
        fl_load_fss     : in     vl_logic;
        fl_load_uds_trn : in     vl_logic;
        fl_erase_cfg0   : in     vl_logic;
        fl_erase_ufm0   : in     vl_logic;
        fl_erase_trim   : in     vl_logic;
        fl_erase_fea    : in     vl_logic;
        fl_load_pkey0   : in     vl_logic;
        fl_load_pkey1   : in     vl_logic;
        fl_load_pkey2   : in     vl_logic;
        fl_load_pkey3   : in     vl_logic;
        fl_load_udss1   : in     vl_logic;
        fl_load_ufs1    : in     vl_logic;
        fl_load_pks     : in     vl_logic;
        fl_load_css     : in     vl_logic;
        fl_load_csec    : in     vl_logic;
        fl_erase_cfg1   : in     vl_logic;
        fl_erase_ufm1   : in     vl_logic;
        fl_erase_pubkey : in     vl_logic;
        fl_erase_csec   : in     vl_logic;
        fl_load_akey0   : in     vl_logic;
        fl_load_akey1   : in     vl_logic;
        fl_load_ufs2    : in     vl_logic;
        fl_load_ufs3    : in     vl_logic;
        fl_load_aks     : in     vl_logic;
        fl_load_uss     : in     vl_logic;
        fl_load_usec    : in     vl_logic;
        fl_erase_ufm2   : in     vl_logic;
        fl_erase_ufm3   : in     vl_logic;
        fl_erase_aeskey : in     vl_logic;
        fl_erase_usec   : in     vl_logic;
        lsc_sdm         : in     vl_logic;
        lsc_sdm_cfg0    : in     vl_logic;
        lsc_sdm_cfg1    : in     vl_logic;
        sdm_start_bse   : in     vl_logic;
        sdm_bse_eof     : in     vl_logic;
        preamble_std_sdm: in     vl_logic;
        preamble_enc_sdm: in     vl_logic;
        preamble_err_sdm: in     vl_logic;
        sram_sec_prog   : in     vl_logic;
        sram_sec_read   : in     vl_logic;
        sram_done       : in     vl_logic;
        sram_ues        : in     vl_logic_vector(31 downto 0);
        sf_exec_buf     : in     vl_logic_vector(127 downto 0);
        busy_sram       : in     vl_logic;
        fail_sram       : in     vl_logic;
        sf_finish_bke   : in     vl_logic;
        fl_exec_buf     : in     vl_logic_vector(127 downto 0);
        fl_modal_state  : in     vl_logic_vector(31 downto 0);
        fl_pg_count     : in     vl_logic_vector(9 downto 0);
        fl_er_count     : in     vl_logic_vector(11 downto 0);
        row             : in     vl_logic_vector(14 downto 6);
        busy_flash      : in     vl_logic;
        fail_flash      : in     vl_logic;
        fail_sdm_a      : in     vl_logic;
        fail_sdm_b      : in     vl_logic;
        fl_busy_ppt     : in     vl_logic;
        fl_busy_cdm     : in     vl_logic;
        fl_busy_sdm     : in     vl_logic;
        fl_finish_ppt   : in     vl_logic;
        fl_finish_cdm   : in     vl_logic;
        fl_finish_sdm   : in     vl_logic;
        ctrl_ndr        : in     vl_logic;
        ctrl_ncdm       : in     vl_logic;
        ctrl_nbke       : in     vl_logic;
        ctrl_ebr_init_en: in     vl_logic;
        ctrl_wkup_tran  : in     vl_logic;
        ctrl_hfc_hd     : in     vl_logic;
        ctrl_mspim_sel  : in     vl_logic;
        ctrl_tran_ebr   : in     vl_logic;
        ctrl_tran_ip    : in     vl_logic;
        ctrl_tran_hse   : in     vl_logic;
        ctrl_tran_edit  : in     vl_logic;
        ctrl_pdone_ovld : in     vl_logic_vector(1 downto 0);
        ctrl_erase_all  : in     vl_logic;
        cib_mspim_addr  : in     vl_logic_vector(15 downto 0);
        cib_mcsn_sel    : in     vl_logic;
        cib_user_gsr    : in     vl_logic;
        cib_tsall       : in     vl_logic;
        mc1_gsr_phase   : in     vl_logic_vector(2 downto 0);
        mc1_gwe_phase   : in     vl_logic_vector(2 downto 0);
        mc1_goe_phase   : in     vl_logic_vector(2 downto 0);
        mc1_done_phase  : in     vl_logic_vector(3 downto 0);
        mc1_pll_chk     : in     vl_logic_vector(7 downto 0);
        mc1_sync_ext_done: in     vl_logic;
        mc1_mspi_sed_addr: in     vl_logic_vector(15 downto 0);
        mc1_source_sel  : in     vl_logic;
        mc1_mspi_addr   : in     vl_logic_vector(15 downto 0);
        mc1_gsrn        : in     vl_logic;
        mc1_goe         : in     vl_logic;
        mc1_gwe         : in     vl_logic;
        mc1_mib         : in     vl_logic;
        mc1_pcs         : in     vl_logic;
        mc1_pupn        : in     vl_logic;
        mc1_en_tsall    : in     vl_logic;
        mc1_tsall_inv   : in     vl_logic;
        mc1_sleep_gsrn  : in     vl_logic;
        mc1_sleep_gwe   : in     vl_logic;
        mc1_sleep_pupn  : in     vl_logic;
        mc1_sleep_fio   : in     vl_logic;
        mc1_gsrn_inv    : in     vl_logic;
        mc1_gsrn_sync   : in     vl_logic;
        mc1_user_gsrn   : in     vl_logic;
        mc1_wkup_pw     : in     vl_logic_vector(3 downto 0);
        mc1_wkup_pd     : in     vl_logic_vector(3 downto 0);
        rti2d           : in     vl_logic;
        rti_r           : in     vl_logic;
        upir_ss_r       : in     vl_logic;
        seldr_ss        : in     vl_logic;
        capdr_ss_r      : in     vl_logic;
        exit1dr_ss_r    : in     vl_logic;
        bsmode1         : in     vl_logic;
        tsall_ctrl      : in     vl_logic;
        isc_enabled     : in     vl_logic;
        isc_disable_completing: in     vl_logic;
        jaccess_sram    : in     vl_logic;
        jaccess_flash   : in     vl_logic;
        jaccess_fl_norm : in     vl_logic;
        jaccess_fl_sudo : in     vl_logic;
        jaccess_fl_safe : in     vl_logic;
        jaccess_tag     : in     vl_logic;
        jaccess_flash_all: in     vl_logic;
        jenable_offl    : in     vl_logic;
        jtag_active     : in     vl_logic;
        j_enable_qual   : in     vl_logic;
        j_enable_x_qual : in     vl_logic;
        jexit_fl_offline: in     vl_logic;
        jexit_normal    : in     vl_logic;
        jexit_fl_tran   : in     vl_logic;
        j_disable_qual  : in     vl_logic;
        jrst_isc_done_i : in     vl_logic;
        jset_isc_done_i : in     vl_logic;
        jconfig_dat     : in     vl_logic_vector(3 downto 0);
        jcontxt_dat     : in     vl_logic_vector(7 downto 0);
        jsector_dat     : in     vl_logic_vector(15 downto 0);
        jbuf128_dat     : in     vl_logic_vector(127 downto 0);
        jburst_en       : in     vl_logic;
        lsc_auth_ctrl_cq: in     vl_logic;
        lsc_verify_uid_cq: in     vl_logic;
        lsc_erase_all_cq: in     vl_logic;
        persist_mspi    : in     vl_logic;
        mc1_erase_all   : in     vl_logic_vector(7 downto 0);
        mfg_en          : in     vl_logic;
        mfg_margin      : in     vl_logic;
        mfg_bkgrndft_en : in     vl_logic;
        mfg_freq_sel    : in     vl_logic;
        isc_data_shift_iq: in     vl_logic;
        isc_addr_shift_iq: in     vl_logic;
        verify_id_iq    : in     vl_logic;
        idcode_pub_iq   : in     vl_logic;
        uidcode_pub_iq  : in     vl_logic;
        usercode_iq     : in     vl_logic;
        usercode_dryrun_iq: in     vl_logic;
        read_temp_iq    : in     vl_logic;
        lsc_device_ctrl_iq: in     vl_logic;
        prog_dryrun_addr_iq: in     vl_logic;
        lsc_shift_password_iq: in     vl_logic;
        lsc_read_status_mq: in     vl_logic;
        lsc_read_status1_iq: in     vl_logic;
        lsc_read_mfg_status_mq: in     vl_logic;
        lsc_refresh_iq  : in     vl_logic;
        lsc_bitstream_burst_iq: in     vl_logic;
        lsc_i2ci_crbr_wt_iq: in     vl_logic;
        lsc_i2ci_txdr_wt_iq: in     vl_logic;
        lsc_i2ci_rxdr_rd_iq: in     vl_logic;
        lsc_i2ci_sr_rd_iq: in     vl_logic;
        idcode_prv_iq   : in     vl_logic;
        lsc_read_pes_mq : in     vl_logic;
        lsc_prog_ctrl0_iq: in     vl_logic;
        lsc_read_ctrl0_iq: in     vl_logic;
        lsc_prog_ctrl1_iq: in     vl_logic;
        lsc_read_ctrl1_iq: in     vl_logic;
        lsc_reset_crc_iq: in     vl_logic;
        lsc_read_crc_iq : in     vl_logic;
        lsc_write_comp_dic_iq: in     vl_logic;
        lsc_read_comp_dic_mq: in     vl_logic;
        sf_prog_ucode_iq: in     vl_logic;
        sf_program_iq   : in     vl_logic;
        sf_read_iq      : in     vl_logic;
        sf_erase_iq     : in     vl_logic;
        sf_prog_done_iq : in     vl_logic;
        sf_erase_done_iq: in     vl_logic;
        sf_prog_sec_iq  : in     vl_logic;
        sf_init_addr_iq : in     vl_logic;
        sf_write_addr_iq: in     vl_logic;
        sf_prog_incr_rti_iq: in     vl_logic;
        sf_prog_incr_enc_iq: in     vl_logic;
        sf_prog_incr_cmp_iq: in     vl_logic;
        sf_prog_incr_cne_iq: in     vl_logic;
        sf_vfy_incr_rti_iq: in     vl_logic;
        sf_prog_sed_crc_iq: in     vl_logic;
        sf_read_sed_crc_iq: in     vl_logic;
        sf_write_bus_addr_iq: in     vl_logic;
        sf_pcs_write_iq : in     vl_logic;
        sf_pcs_read_iq  : in     vl_logic;
        sf_ebr_write_iq : in     vl_logic;
        sf_ebr_read_iq  : in     vl_logic;
        fl_prog_ucode_iq: in     vl_logic;
        fl_erase_iq     : in     vl_logic;
        fl_prog_done_iq : in     vl_logic;
        fl_prog_sec_iq  : in     vl_logic;
        fl_prog_secplus_iq: in     vl_logic;
        fl_init_addr_iq : in     vl_logic;
        fl_write_addr_iq: in     vl_logic;
        fl_prog_incr_nv_iq: in     vl_logic;
        fl_read_incr_nv_iq: in     vl_logic;
        fl_prog_password_iq: in     vl_logic;
        fl_read_password_iq: in     vl_logic;
        fl_prog_cipher_key0_iq: in     vl_logic;
        fl_read_cipher_key0_iq: in     vl_logic;
        fl_prog_cipher_key1_iq: in     vl_logic;
        fl_read_cipher_key1_iq: in     vl_logic;
        fl_prog_feature_iq: in     vl_logic;
        fl_read_feature_iq: in     vl_logic;
        fl_prog_feabits_iq: in     vl_logic;
        fl_read_feabits_iq: in     vl_logic;
        fl_init_addr_ufm_iq: in     vl_logic;
        fl_prog_tag_iq  : in     vl_logic;
        fl_erase_tag_iq : in     vl_logic;
        fl_read_tag_iq  : in     vl_logic;
        fl_prog_pes_mq  : in     vl_logic;
        fl_prog_trim0_mq: in     vl_logic;
        fl_prog_trim1_mq: in     vl_logic;
        fl_prog_mes_mq  : in     vl_logic;
        fl_prog_hes_mq  : in     vl_logic;
        fl_read_trim0_mq: in     vl_logic;
        fl_read_trim1_mq: in     vl_logic;
        fl_read_mes_mq  : in     vl_logic;
        fl_read_hes_mq  : in     vl_logic;
        fl_prog_csec_iq : in     vl_logic;
        fl_read_csec_iq : in     vl_logic;
        fl_prog_usec_iq : in     vl_logic;
        fl_read_usec_iq : in     vl_logic;
        fl_prog_authdone_iq: in     vl_logic;
        fl_prog_authmode_iq: in     vl_logic;
        fl_prog_aesfea_iq: in     vl_logic;
        fl_read_authmode_iq: in     vl_logic;
        fl_read_aesfea_iq: in     vl_logic;
        mfg_mtest_mq    : in     vl_logic;
        mfg_mtrim_mq    : in     vl_logic;
        mfg_mdata_mq    : in     vl_logic;
        mfg_bist_status_mq: in     vl_logic;
        mfg_bist_en_mq  : in     vl_logic;
        mem_bist_status : in     vl_logic_vector(127 downto 0);
        isc_nj_enabled  : in     vl_logic;
        isc_nj_disable_completing: in     vl_logic;
        njaccess_sram   : in     vl_logic;
        njaccess_flash  : in     vl_logic;
        njaccess_fl_norm: in     vl_logic;
        njaccess_fl_sudo: in     vl_logic;
        njaccess_fl_safe: in     vl_logic;
        njaccess_tag    : in     vl_logic;
        njaccess_flash_all: in     vl_logic;
        njenable_offl   : in     vl_logic;
        njtag_active    : in     vl_logic;
        njtag_active_nsed: in     vl_logic;
        nj_enable_qual  : in     vl_logic;
        nj_enable_x_qual: in     vl_logic;
        nj_exec_a       : in     vl_logic;
        nj_exec_b       : in     vl_logic;
        nj_exec_c       : in     vl_logic;
        nj_exec_d       : in     vl_logic;
        nj_exec_e       : in     vl_logic;
        nj_exec_f       : in     vl_logic;
        njexit_fl_offline: in     vl_logic;
        njexit_normal   : in     vl_logic;
        njexit_fl_tran  : in     vl_logic;
        nj_disable_qual : in     vl_logic;
        njrst_isc_done_c: in     vl_logic;
        njset_isc_done_c: in     vl_logic;
        njconfig_dat    : in     vl_logic_vector(3 downto 0);
        njcontxt_dat    : in     vl_logic_vector(7 downto 0);
        njsector_dat    : in     vl_logic_vector(15 downto 0);
        njbuf128_dat    : in     vl_logic_vector(127 downto 0);
        bse_end_cqual   : in     vl_logic;
        njm_invalid_c   : in     vl_logic;
        njr_invalid_c   : in     vl_logic;
        njs_invalid_c   : in     vl_logic;
        sed_invalid_c   : in     vl_logic;
        nj_jump_param   : in     vl_logic_vector(31 downto 0);
        nj_csel_param   : in     vl_logic_vector(7 downto 0);
        njburst_inp     : in     vl_logic;
        isc_data_shift_cq: in     vl_logic;
        isc_addr_shift_cq: in     vl_logic;
        verify_id_cq    : in     vl_logic;
        idcode_pub_cq   : in     vl_logic;
        uidcode_pub_cq  : in     vl_logic;
        usercode_cq     : in     vl_logic;
        usercode_dryrun_cq: in     vl_logic;
        read_temp_cq    : in     vl_logic;
        lsc_device_ctrl_cq: in     vl_logic;
        prog_dryrun_addr_cq: in     vl_logic;
        lsc_shift_password_cq: in     vl_logic;
        lsc_read_status_cq: in     vl_logic;
        lsc_read_status1_cq: in     vl_logic;
        lsc_check_busy_cq: in     vl_logic;
        lsc_refresh_cq  : in     vl_logic;
        lsc_bitstream_burst_cq: in     vl_logic;
        lsc_i2ci_crbr_wt_cq: in     vl_logic;
        lsc_i2ci_txdr_wt_cq: in     vl_logic;
        lsc_i2ci_rxdr_rd_cq: in     vl_logic;
        lsc_i2ci_sr_rd_cq: in     vl_logic;
        idcode_prv_cq   : in     vl_logic;
        lsc_read_pes_cq : in     vl_logic;
        lsc_prog_ctrl0_cq: in     vl_logic;
        lsc_read_ctrl0_cq: in     vl_logic;
        lsc_prog_ctrl1_cq: in     vl_logic;
        lsc_read_ctrl1_cq: in     vl_logic;
        lsc_reset_crc_cq: in     vl_logic;
        lsc_read_crc_cq : in     vl_logic;
        lsc_write_comp_dic_cq: in     vl_logic;
        sf_prog_ucode_cq: in     vl_logic;
        sf_program_cq   : in     vl_logic;
        sf_read_cq      : in     vl_logic;
        sf_erase_cq     : in     vl_logic;
        sf_prog_done_cq : in     vl_logic;
        sf_erase_done_cq: in     vl_logic;
        sf_prog_sec_cq  : in     vl_logic;
        sf_init_addr_cq : in     vl_logic;
        sf_write_addr_cq: in     vl_logic;
        sf_prog_incr_rti_cq: in     vl_logic;
        sf_prog_incr_enc_cq: in     vl_logic;
        sf_prog_incr_cmp_cq: in     vl_logic;
        sf_prog_incr_cne_cq: in     vl_logic;
        sf_vfy_incr_rti_cq: in     vl_logic;
        sf_prog_sed_crc_cq: in     vl_logic;
        sf_read_sed_crc_cq: in     vl_logic;
        sf_write_bus_addr_cq: in     vl_logic;
        sf_pcs_write_cq : in     vl_logic;
        sf_pcs_read_cq  : in     vl_logic;
        sf_ebr_write_cq : in     vl_logic;
        sf_ebr_read_cq  : in     vl_logic;
        fl_prog_ucode_cq: in     vl_logic;
        fl_erase_cq     : in     vl_logic;
        fl_prog_done_cq : in     vl_logic;
        fl_prog_sec_cq  : in     vl_logic;
        fl_prog_secplus_cq: in     vl_logic;
        fl_init_addr_cq : in     vl_logic;
        fl_write_addr_cq: in     vl_logic;
        fl_prog_incr_nv_cq: in     vl_logic;
        fl_read_incr_nv_cq: in     vl_logic;
        fl_prog_password_cq: in     vl_logic;
        fl_read_password_cq: in     vl_logic;
        fl_prog_cipher_key0_cq: in     vl_logic;
        fl_read_cipher_key0_cq: in     vl_logic;
        fl_prog_cipher_key1_cq: in     vl_logic;
        fl_read_cipher_key1_cq: in     vl_logic;
        fl_prog_feature_cq: in     vl_logic;
        fl_read_feature_cq: in     vl_logic;
        fl_prog_feabits_cq: in     vl_logic;
        fl_read_feabits_cq: in     vl_logic;
        fl_init_addr_ufm_cq: in     vl_logic;
        fl_prog_tag_cq  : in     vl_logic;
        fl_erase_tag_cq : in     vl_logic;
        fl_read_tag_cq  : in     vl_logic;
        fl_prog_csec_cq : in     vl_logic;
        fl_read_csec_cq : in     vl_logic;
        fl_prog_usec_cq : in     vl_logic;
        fl_read_usec_cq : in     vl_logic;
        fl_prog_authdone_cq: in     vl_logic;
        fl_prog_authmode_cq: in     vl_logic;
        fl_prog_aesfea_cq: in     vl_logic;
        fl_read_authmode_cq: in     vl_logic;
        fl_read_aesfea_cq: in     vl_logic;
        lsc_jump_cq     : in     vl_logic;
        lsc_chip_select_cq: in     vl_logic;
        lsc_flow_through_cq: in     vl_logic;
        bypass_cq       : in     vl_logic;
        sed_init_addr_cq: in     vl_logic;
        sed_write_addr_cq: in     vl_logic;
        sed_prog_incr_rti_cq: in     vl_logic;
        sed_prog_incr_cmp_cq: in     vl_logic;
        sed_prog_sed_crc_cq: in     vl_logic;
        sed_prog_ctrl0_cq: in     vl_logic;
        sed_prog_ctrl1_cq: in     vl_logic;
        sed_write_comp_dic_cq: in     vl_logic;
        cib_pll_lock    : in     vl_logic_vector(7 downto 0);
        sf_asr_out      : in     vl_logic;
        fl_prog_pubkey0_cq: in     vl_logic;
        fl_read_pubkey0_cq: in     vl_logic;
        fl_prog_pubkey0_iq: in     vl_logic;
        fl_read_pubkey0_iq: in     vl_logic;
        fl_prog_pubkey1_cq: in     vl_logic;
        fl_read_pubkey1_cq: in     vl_logic;
        fl_prog_pubkey1_iq: in     vl_logic;
        fl_read_pubkey1_iq: in     vl_logic;
        fl_prog_pubkey2_cq: in     vl_logic;
        fl_read_pubkey2_cq: in     vl_logic;
        fl_prog_pubkey2_iq: in     vl_logic;
        fl_read_pubkey2_iq: in     vl_logic;
        fl_prog_pubkey3_cq: in     vl_logic;
        fl_read_pubkey3_cq: in     vl_logic;
        fl_prog_pubkey3_iq: in     vl_logic;
        fl_read_pubkey3_iq: in     vl_logic;
        key_rst_sync    : in     vl_logic;
        key_shift_en    : in     vl_logic;
        lsc_alter_sec_cq: in     vl_logic;
        lsc_alter_sram_sec_cq: in     vl_logic;
        lsc_alter_port_sec_cq: in     vl_logic;
        lsc_prog_uds_cq : in     vl_logic;
        p_iboot0s       : in     vl_logic;
        dec_ready       : in     vl_logic;
        auth_en         : in     vl_logic;
        auth_ready      : in     vl_logic;
        auth_fail       : in     vl_logic;
        auth_done       : in     vl_logic;
        auth_time_out   : in     vl_logic;
        auth_setup_fail : in     vl_logic;
        auth_bs_err     : in     vl_logic;
        tc_to           : in     vl_logic;
        tc_to_reboot_en : in     vl_logic;
        tc_to_reboot_mode: in     vl_logic;
        isc_prog_done_c : in     vl_logic;
        hse_trn_dat     : in     vl_logic_vector(127 downto 0);
        cib_thr_det_clk : in     vl_logic;
        cib_thr_det_en  : in     vl_logic;
        cib_lck_thr_src : in     vl_logic;
        mc1_port_lock_en: in     vl_logic_vector(1 downto 0);
        cib_thr_det     : out    vl_logic;
        cib_thr_typ     : out    vl_logic_vector(1 downto 0);
        cib_thr_src     : out    vl_logic_vector(1 downto 0);
        passwordThrDetEnable: in     vl_logic;
        accessLockSectorDetEnable: in     vl_logic;
        illegalManuModeDetEnable: in     vl_logic;
        JTAGThrDetEnable: in     vl_logic;
        slaveSPIThrDetEnable: in     vl_logic;
        slaveI2CThrDetEnable: in     vl_logic;
        wishboneThrDetEnable: in     vl_logic;
        jsel_mfg        : in     vl_logic;
        sspi_active     : in     vl_logic;
        i2c_active      : in     vl_logic
    );
end cfg_cntl;
