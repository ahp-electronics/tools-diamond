library verilog;
use verilog.vl_types.all;
entity hse_top_wrap is
    port(
        por_n           : in     vl_logic;
        clk_osc         : in     vl_logic;
        reset           : in     vl_logic;
        scan_mode       : in     vl_logic;
        enc_enabled     : in     vl_logic;
        wb_clk_i        : in     vl_logic;
        wb_rst_i        : in     vl_logic;
        wb_stb_i        : in     vl_logic;
        wb_cyc_i        : in     vl_logic;
        wb_we_i         : in     vl_logic;
        wb_dat_i        : in     vl_logic_vector(31 downto 0);
        wb_adr_i        : in     vl_logic_vector(17 downto 0);
        wb_dat_o        : out    vl_logic_vector(31 downto 0);
        wb_ack_o        : out    vl_logic;
        asf_reset_i     : in     vl_logic;
        asf_clk_i       : in     vl_logic;
        asf_wr_i        : in     vl_logic;
        asf_full_o      : out    vl_logic;
        asf_empty_o     : out    vl_logic;
        asf_rd_i        : in     vl_logic;
        cfg_clk         : in     vl_logic;
        off_hse_usrmd   : in     vl_logic;
        cfg_active      : in     vl_logic;
        cfg_noise       : in     vl_logic;
        ac_alg_sel      : in     vl_logic_vector(1 downto 0);
        data_in         : in     vl_logic_vector(7 downto 0);
        write_en        : in     vl_logic;
        last_cbyte      : in     vl_logic;
        busy            : out    vl_logic_vector(1 downto 0);
        buffer_ready    : out    vl_logic;
        pass_fail       : out    vl_logic;
        pf_valid        : out    vl_logic;
        uds_out         : out    vl_logic_vector(255 downto 0);
        uds_in          : in     vl_logic_vector(255 downto 0);
        ebr_hse_spram_0_BistFail: out    vl_logic;
        ebr_hse_spram_0_ErrMap: out    vl_logic;
        ebr_hse_spram_0_Finish: out    vl_logic;
        ebr_hse_spram_0_BistEn: in     vl_logic;
        ebr_hse_spram_1_BistFail: out    vl_logic;
        ebr_hse_spram_1_ErrMap: out    vl_logic;
        ebr_hse_spram_1_Finish: out    vl_logic;
        ebr_hse_spram_1_BistEn: in     vl_logic;
        ebr_hse_spram_2_BistFail: out    vl_logic;
        ebr_hse_spram_2_ErrMap: out    vl_logic;
        ebr_hse_spram_2_Finish: out    vl_logic;
        ebr_hse_spram_2_BistEn: in     vl_logic;
        ebr_hse_spram_3_BistFail: out    vl_logic;
        ebr_hse_spram_3_ErrMap: out    vl_logic;
        ebr_hse_spram_3_Finish: out    vl_logic;
        ebr_hse_spram_3_BistEn: in     vl_logic;
        ebr_hse_spram_4_BistFail: out    vl_logic;
        ebr_hse_spram_4_ErrMap: out    vl_logic;
        ebr_hse_spram_4_Finish: out    vl_logic;
        ebr_hse_spram_4_BistEn: in     vl_logic;
        ebr_hse_spram_5_BistFail: out    vl_logic;
        ebr_hse_spram_5_ErrMap: out    vl_logic;
        ebr_hse_spram_5_Finish: out    vl_logic;
        ebr_hse_spram_5_BistEn: in     vl_logic;
        ebr_hse_spram_6_BistFail: out    vl_logic;
        ebr_hse_spram_6_ErrMap: out    vl_logic;
        ebr_hse_spram_6_Finish: out    vl_logic;
        ebr_hse_spram_6_BistEn: in     vl_logic;
        ebr_hse_spram_7_BistFail: out    vl_logic;
        ebr_hse_spram_7_ErrMap: out    vl_logic;
        ebr_hse_spram_7_Finish: out    vl_logic;
        ebr_hse_spram_7_BistEn: in     vl_logic;
        ebr_hse_Bisted_rom64kx32_BistFail: out    vl_logic;
        ebr_hse_Bisted_rom64kx32_SignatureParallel: out    vl_logic_vector(49 downto 0);
        ebr_hse_Bisted_rom64kx32_Finsh: out    vl_logic;
        ebr_hse_Bisted_rom64kx32_BistEn: in     vl_logic;
        ebr_hse_Bisted_rom4kx32_BistFail: out    vl_logic;
        ebr_hse_Bisted_rom4kx32_SignatureParallel: out    vl_logic_vector(49 downto 0);
        ebr_hse_Bisted_rom4kx32_Finsh: out    vl_logic;
        ebr_hse_Bisted_rom4kx32_BistEn: in     vl_logic
    );
end hse_top_wrap;
