library verilog;
use verilog.vl_types.all;
entity pcs_quad_clk_mux is
    port(
        sysclk0         : out    vl_logic;
        sysclk1         : out    vl_logic;
        sysclk2         : out    vl_logic;
        sysclk3         : out    vl_logic;
        pcs_rxclk0      : out    vl_logic;
        pcs_rxclk1      : out    vl_logic;
        pcs_rxclk2      : out    vl_logic;
        pcs_rxclk3      : out    vl_logic;
        m_rxclk0        : out    vl_logic;
        m_rxclk1        : out    vl_logic;
        m_rxclk2        : out    vl_logic;
        m_rxclk3        : out    vl_logic;
        fb_rxclk0       : out    vl_logic;
        fb_rxclk1       : out    vl_logic;
        fb_rxclk2       : out    vl_logic;
        fb_rxclk3       : out    vl_logic;
        sysclk0_slow    : out    vl_logic;
        sysclk1_slow    : out    vl_logic;
        sysclk2_slow    : out    vl_logic;
        sysclk3_slow    : out    vl_logic;
        fb_rxclk0_slow  : out    vl_logic;
        fb_rxclk1_slow  : out    vl_logic;
        fb_rxclk2_slow  : out    vl_logic;
        fb_rxclk3_slow  : out    vl_logic;
        txclk0          : in     vl_logic;
        txclk1          : in     vl_logic;
        txclk2          : in     vl_logic;
        txclk3          : in     vl_logic;
        rxclk0          : in     vl_logic;
        rxclk1          : in     vl_logic;
        rxclk2          : in     vl_logic;
        rxclk3          : in     vl_logic;
        cascade_clk     : in     vl_logic;
        test_clk        : in     vl_logic;
        pcs_mode        : in     vl_logic;
        uc_mode         : in     vl_logic;
        x4_mode         : in     vl_logic;
        cascade_en      : in     vl_logic;
        mclksel_0       : in     vl_logic_vector(1 downto 0);
        mclksel_1       : in     vl_logic_vector(1 downto 0);
        mclksel_2       : in     vl_logic_vector(1 downto 0);
        mclksel_3       : in     vl_logic_vector(1 downto 0);
        sb_loopback_0   : in     vl_logic;
        sb_loopback_1   : in     vl_logic;
        sb_loopback_2   : in     vl_logic;
        sb_loopback_3   : in     vl_logic;
        scan_mode       : in     vl_logic;
        test_mode       : in     vl_logic_vector(2 downto 0)
    );
end pcs_quad_clk_mux;
