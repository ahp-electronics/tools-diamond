library verilog;
use verilog.vl_types.all;
entity vlov1mce is
    port(
        Z               : out    vl_logic
    );
end vlov1mce;
