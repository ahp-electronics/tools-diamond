library verilog;
use verilog.vl_types.all;
entity oa_22222222 is
    port(
        A               : in     vl_logic_vector(7 downto 0);
        EN              : in     vl_logic_vector(7 downto 0);
        Z               : out    vl_logic
    );
end oa_22222222;
