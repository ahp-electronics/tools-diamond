--
@ER--B$FbsEHo0OR52gR4g-cRRj.jd$R1MHbDO$H0ROQM
R--fN]C8:CsR#//$DMbH0OH$N/lb..jjDjdNl0/NCbbsN#/0D0/HoL/CFM_s.ONNN/sl__sIE3P8Ry4f-
-
-

--
-Rl1HbRDC)RqvIEH0Rb#CC0sNC7Rq71) 1FRVsCRsNN8RMI8RsCH0
R--aoNsC:0RROpkCRM0-)RmB.qRq-
-

--
LDHs$NsRCHCCk;
#HCRC3CC#_08DHFoO4_4nNc3D
D;kR#CHCCC38#0_oDFH#O_HCoM8D3NDD;
HNLssF$Rs.ON;#
kCsRFO3N.FNsOObFl3DND;M
C0$H0Rv)q_W)_R
H#RRRRoCCMsRHO5R
RRRRRRNRVl$HD:0R#soHMRR:="MMFC
";RRRRRRRRI0H8ERR:HCM0oRCs:4=R;RR
RRRRRNRR8I8sHE80RH:RMo0CC:sR=;RcRRRRRRRR-L-RHCoRMoFkEFRVsCR8b
0ERRRRRRRR80CbERR:HCM0oRCs:R=R4
n;RRRRRRRR80Fk_osCRL:RFCFDN:MR=NRVD;#CRRRRRR--ERN#Fbk0ks0RCRo
RRRRR8RRHsM_C:oRRFLFDMCNRR:=V#NDCR;RRRRR-E-RN8#RNR0NHkMb0CRsoR
RRRRRRNRs8_8ssRCo:FRLFNDCM=R:RDVN#RC;R-RR-NRE8CRsNN8R8C8s#s#RCRo
RRRRRIRRNs88_osCRL:RFCFDN:MR=NRVDR#CRRRR-E-RNI8RsCH0R8N8s#C#RosC
RRRRRRRR
2;RRRRb0FsRR5
RRRRR7RRmRzaRF:Rk#0R0D8_FOoH_OPC05FsI0H8ER-48MFI0jFR2R;
RRRRR)RRq)77RH:RM#RR0D8_FOoH_OPC05FsNs88I0H8ER-48MFI0jFR2R;
RRRRR7RRQRhRRH:RM#RR0D8_FOoH_OPC05FsI0H8ER-48MFI0jFR2R;
RRRRRWRRq)77RH:RM#RR0D8_FOoH_OPC05FsNs88I0H8ER-48MFI0jFR2R;
RRRRRWRR RRRRH:RM#RR0D8_FOoH;RRRRRRR-I-RsCH0RNCMLRDCVRFss
NlRRRRRRRRBRpiRRR:HRMR#_08DHFoOR;RRRRRRR--OODF	FRVsNRslN,R8,8sRM8H
RRRRRRRRpmBi:RRRRHMR8#0_oDFHRORRRRRR-R-R0FbRFODOV	RF8sRF
k0RRRRRRRR2C;
MC8RM00H$qR)v__)W
;
---
-HRwsR#0HDlbCMlC0HN0FlMRkR#0LOCRNCDD8sRNO
Ej-N-
sHOE00COkRsCNEsOjVRFRv)q_W)_R
H#O#FM00NMRlMk_DOCD8#_CRCb:MRH0CCos=R:R855CEb0R4-R2n/42R;RRRRRR-RR-RRyFsVRFRI#F7VRBnw4XR.ZODCD#CRMC88C
MOF#M0N0kRMlC_OD_D#ICH8RH:RMo0CC:sR=5R5I0H8ERR-4.2/2R;RRRRRRRRR-y-RRRFVOkFDlRM#F7VRBnw4XR.ZODCD#CRMC88C
o#HMRNDF_k0CRMRRRR:#_08DHFoOC_POs0F5lMk_DOCD8#_CRCb8MFI0jFR2R;R-C-RMDNLCV#RF0sRs#H-0CN0#H
#oDMNRCIb_RCMR:RRR8#0_oDFHPO_CFO0sk5MlC_OD_D#8bCCRI8FMR0FjR2;RR--I0sHCMRCNCLD#FRVsNRCOsERFFIRVqR)vCROD
D##MHoNHDRMC_soRRRR#:R0D8_FOoH_OPC05FsI0H8ER+48MFI0jFR2R;RRRRRR-RR-#RkC08RFCRso0H#C7sRQ
hR#MHoNFDRks0_CRoRR#:R0D8_FOoH_OPC05FsI0H8ER+48MFI0jFR2R;RRRRRR-RR-#RkC08RFCRso0H#C7sRm
za#MHoNsDRNs8_CRoRR#:R0D8_FOoH_OPC05FsNs88I0H8ER-48MFI0jFR2R;RR-RR-#RkC08RFCRso0H#C)sRq)77
o#HMRNDI_N8sRCoRRR:#_08DHFoOC_POs0F58N8s8IH04E-RI8FMR0FjR2;RRRR-k-R#RC80sFRC#oH0RCsW7q7)H
#oDMNRIDF_8sN8:sRR8#0_oDFHPO_CFO0sR5d8MFI0jFR2R;RRRRRRRRRRRRRRR--s8N8sHRL0H#RM0bkRR0F)RqvODCD#cR5R0LH#CRsJskHC
82#MHoNDDRFII_Ns88R#:R0D8_FOoH_OPC05FsdFR8IFM0R;j2RRRRRRRRRRRRR-RR-NRI8R8sL#H0RbHMk00RFqR)vCRODRD#5LcRHR0#skCJH8sC2L

CMoH
R
RR-R-RRQVNs88I0H8ERR<c#RN#MHoR''jRR0Fk#MkCL8RH
0#RRRRzR4R:VRHR85N8HsI8R0E=2R4RMoCC0sNCR
RRRRRRFRDIN_s8R8s<"=Rj"jjRs&RNs8_Cjo52R;
RRRRRDRRFII_Ns88RR<="jjj"RR&I_N8s5Coj
2;RRRRCRM8oCCMsCN0R;z4
RRRRRz.RH:RVNR58I8sHE80R.=R2CRoMNCs0RC
RRRRRDRRFsI_Ns88RR<=""jjRs&RNs8_C4o5RI8FMR0Fj
2;RRRRRRRRD_FII8N8s=R<Rj"j"RR&I_N8s5Co4FR8IFM0R;j2
RRRR8CMRMoCC0sNC.Rz;R
RRdRzRRR:H5VRNs88I0H8ERR=do2RCsMCN
0CRRRRRRRRD_FIs8N8s=R<R''jRs&RNs8_C.o5RI8FMR0Fj
2;RRRRRRRRD_FII8N8s=R<R''jRI&RNs8_C.o5RI8FMR0Fj
2;RRRRCRM8oCCMsCN0R;zd
RRRRRzcRH:RVNR58I8sHE80Rd>R2CRoMNCs0RC
RRRRRDRRFsI_Ns88RR<=s_N8s5CodFR8IFM0R;j2
RRRRRRRRIDF_8IN8<sR=NRI8C_soR5d8MFI0jFR2R;
RCRRMo8RCsMCNR0Cz
c;
RRRRR--Q5VR8_HMs2CoRosCHC#0sQR7h#RkHRMoB
piRRRRzR6R:VRHRH58MC_soo2RCsMCN
0CRRRRRRRRbOsFCR##5iBp,QR7hL2RCMoH
RRRRRRRRRRRRRHV5iBpR'=R4N'RMB8RpCi'P0CM2ER0CRM
RRRRRRRRRRRRRHRRMC_so=R<Rj5"j&"RRh7Q2R;
RRRRRRRRRCRRMH8RVR;
RRRRRCRRMb8RsCFO#
#;RRRRCRM8oCCMsCN0R;z6
RRRRRznRH:RVMR5F80RHsM_CRo2oCCMsCN0
RRRRRRRRRRRR_HMsRCo<5=R""jjR7&RQ;h2
RRRR8CMRMoCC0sNCnRz;R

R-RR-VRQRF58ks0_CRo2sHCo#s0CRz7ma#RkHRMomiBp
RRRRRz(RH:RV8R5F_k0s2CoRMoCC0sNCR
RRRRRRsRbF#OC#mR5B,piR0Fk_osC2CRLo
HMRRRRRRRRRRRRH5VRmiBpR'=R4N'RMm8RB'piCMPC002RE
CMRRRRRRRRRRRRRRRR7amzRR<=F_k0s5CoI0H8ER-48MFI0jFR2R;
RRRRRRRRRCRRMH8RVR;
RRRRRCRRMb8RsCFO#
#;RRRRRRRRCRM8oCCMsCN0R;z(
RRRRRzURH:RVMR5F80RF_k0s2CoRMoCC0sNCR
RRRRRRRRRRmR7z<aR=kRF0C_soH5I8-0E4FR8IFM0R;j2
RRRR8CMRMoCC0sNCURz;R

R-RR-VRQRN5s8_8ss2CoRosCHC#0sqR)7R7)kM#HopRBiR
RRgRzRRR:H5VRs8N8sC_soo2RCsMCN
0CRRRRRRRRbOsFCR##5pmBi),Rq)772CRLo
HMRRRRRRRRRRRRH5VRmiBpR'=R4N'RMm8RB'piCMPC002RE
CMRRRRRRRRRRRRRRRRs_N8sRCo<)=Rq)7758N8s8IH04E-RI8FMR0Fj
2;RRRRRRRRRRRRCRM8H
V;RRRRRRRRCRM8bOsFC;##
RRRR8CMRMoCC0sNCgRz;R
RR4RzjRR:H5VRMRF0s8N8sC_soo2RCsMCN
0CRRRRRRRRRRRRs_N8sRCo<)=Rq)77;R
RRMRC8CRoMNCs0zCR4
j;RRRRRRRR
RRRRR--Q5VRI8N8sC_sos2RC#oH0RCsW7q7)#RkHRMoB
piRRRRzR46RH:RVIR5Ns88_osC2CRoMNCs0RC
RRRRRbRRsCFO#5#RB,piR7Wq7R)2LHCoMR
RRRRRRRRRRVRHRp5BiRR='R4'NRM8B'piCMPC002RE
CMRRRRRRRRRRRRRRRRI_N8sRCo<W=Rq)7758N8s8IH04E-RI8FMR0Fj
2;RRRRRRRRRRRRCRM8H
V;RRRRRRRRCRM8bOsFC;##
RRRR8CMRMoCC0sNC4Rz6R;
RzRR4:nRRRHV50MFR8IN8ss_CRo2oCCMsCN0
RRRRRRRRRRRR8IN_osCRR<=W7q7)R;
RCRRMo8RCsMCNR0Cz;4n
R
RR-R-RMtCC0sNCER0CqR)vCRODRD#NRM8#CCDOD0RFOoH
RRRR4z4RV:RFHsRRRHMM_klODCD#C_8C8bRF0IMFRRjoCCMsCN0
RRRRR--Q5VRNs88I0H8ERR>cM2RCRC80OFRs0CNCsRIHR0CCLMNDNCRMF8Rkk0b0MRCNCLDRD#CCRO0DHFoOR
RRRRRR4Rz.RR:H5VRNs88I0H8ERR>co2RCsMCN
0CRRRRRRRRRRRRRRRRF_k0CHM52=R<R''jRCIEMsR5Ns8_CNo58I8sHE80-84RF0IMF2RcRH=R2DRC#'CR4
';RRRRRRRRRRRRRRRRI_bCCHM52=R<R''4RCIEMIR5Ns8_CNo58I8sHE80-84RF0IMF2RcRH=R2DRC#'CRj
';RRRRRRRRRRRRCRM8oCCMsCN0R.z4;R
RR-R-RRQV58N8s8IH0<ER=2RcRRMFI0sHCMRCNCLDRRFsFbk0kC0RMDNLCCR#D0CORoDFHMORCCC88R
RR4RzdRR:H5VRNs88I0H8E=R<RRc2oCCMsCN0
RRRRRRRRRRRR0Fk_5CMH<2R=jR''R;
RRRRRRRRRRRRRIRRbCC_M25HRR<=';4'
RRRRRRRRRRRR8CMRMoCC0sNC4RzdR;
R-RR-MRtC0sNCER0CqR)vCRODRD#IEH0RH0s-N#00
C#RRRRRRRRzR4c:FRVsRR[HMMRkOl_C#DD_8IHCFR8IFM0RojRCsMCN
0CRRRRRRRRRRRRzv)q:BR7wX4n.
ZRRRRRRRRRRRRRb0FsRblNR)5aQ>R=R0Fk_5CMHR2,7RQj=H>RMC_so.55*2[2,QR74>R=R_HMs5Co5[.*22+4,RR
RRRRRRRRRRRRRRRRRRRRRRRRRjq7RR=>D_FII8N8s25j,7Rq4>R=RIDF_8IN84s52q,R7=.R>FRDIN_I858s.R2,qR7d=D>RFII_Ns885,d2
RRRRRRRRRRRRRRRRRRRRRRRR)RRqR7j=D>RFsI_Ns885,j2R7)q4>R=RIDF_8sN84s52),RqR7.=D>RFsI_Ns885,.2R7)qd>R=RIDF_8sN8ds52R,
RRRRRRRRRRRRRRRRRRRRRRRRR W)h>R=R,W R WuRR=>I_bCCHM52B,Ri>R=RiBp,7R)m=jR>kRF0C_so[55*2.2,7R)m=4R>kRF0C_so[55*+.24;22
RRRRRRRRRRRR8CMRMoCC0sNC4RzcR;
RRRRRCRRMo8RCsMCNR0Cz;44
RRRRRRRRRRRRRRRRRRRRRRRRRRRRCR
MN8RsHOE00COkRsCNEsOj
;

