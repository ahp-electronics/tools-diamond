library verilog;
use verilog.vl_types.all;
entity pcs_mca_control is
    port(
        mrxclk_0        : in     vl_logic;
        mrxclk_2        : in     vl_logic;
        mrxrst0_n       : in     vl_logic;
        mrxrst2_n       : in     vl_logic;
        sync_status_0   : in     vl_logic;
        sync_status_1   : in     vl_logic;
        sync_status_2   : in     vl_logic;
        sync_status_3   : in     vl_logic;
        oof_status_0    : in     vl_logic;
        oof_status_1    : in     vl_logic;
        oof_status_2    : in     vl_logic;
        oof_status_3    : in     vl_logic;
        data_i_0        : in     vl_logic_vector(10 downto 0);
        data_i_1        : in     vl_logic_vector(10 downto 0);
        data_i_2        : in     vl_logic_vector(10 downto 0);
        data_i_3        : in     vl_logic_vector(10 downto 0);
        pcs_mode        : in     vl_logic;
        uc_mode         : in     vl_logic;
        x4_mode         : in     vl_logic;
        x2_mode         : in     vl_logic_vector(1 downto 0);
        rio_mode        : in     vl_logic;
        udf_align_mask  : in     vl_logic_vector(9 downto 0);
        udf_align_a     : in     vl_logic_vector(9 downto 0);
        udf_align_b     : in     vl_logic_vector(9 downto 0);
        mca_ap_0        : in     vl_logic;
        mca_ap_1        : in     vl_logic;
        mca_ap_2        : in     vl_logic;
        mca_ap_3        : in     vl_logic;
        align_en        : in     vl_logic_vector(3 downto 0);
        ab_aligned      : in     vl_logic;
        cd_aligned      : in     vl_logic;
        ab_failed       : in     vl_logic;
        cd_failed       : in     vl_logic;
        asm_disable_ab  : in     vl_logic;
        asm_disable_cd  : in     vl_logic;
        sm_reset_ab_n   : out    vl_logic;
        sm_reset_cd_n   : out    vl_logic;
        pp_ap_0         : out    vl_logic;
        pp_ap_1         : out    vl_logic;
        pp_ap_2         : out    vl_logic;
        pp_ap_3         : out    vl_logic;
        align_status_ab : out    vl_logic;
        align_status_cd : out    vl_logic;
        cascade_en      : in     vl_logic;
        cascade_and_fp  : in     vl_logic;
        cascade_or_fp   : in     vl_logic;
        quad_and_fp_bus : out    vl_logic_vector(1 downto 0);
        quad_or_fp_bus  : out    vl_logic_vector(1 downto 0)
    );
end pcs_mca_control;
