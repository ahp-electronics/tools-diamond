--
@ER--RbBF$osHE50RO42RgRgg1b$MDHHO0R$,Q3MO
R--RDqDRosHER0#sCC#s8PC3-
-
R--#CCDOF0HMCR#0CR8VHHM0MHF3WRRCHRIDCDRP0CMkDND$8RN8DRLF_O	sRFl0
FF-N-RsDOEHR#0=CR#D0CO_lsF

---f-R]8CNCRs:/$/#MHbDO$H0/blN.jj.jNdD0N/lbsbC#H/GDGHM/LDH/MoCCOsH/MoC_MoCCOsH/lsF38PEyf4R

--
LDHs$NsRCHCC
;
kR#CHCCC38#0_oDFH4O_43ncN;DD
Ck#RCHCC03#8F_Do_HON0sHED3NDk;
#HCRC3CC#_08DHFoOM_k#MHoCN83D
D;kR#CI	Fs3MoCb	NON3oCN;DD
H
DLssN$MRkHl#H;#
kCMRkHl#H3FPOlMbFC#M03DND;C

M00H$mR)vN_L#HCR#o
SCsMCH5OR
SSSI0H8ERR:HCM0oRCs:c=R;S
SS8N8s8IH0:ERR0HMCsoCRR:=(S;
SFSDI8N8sRR:HCM0oRCs:j=R;S
SSoEHE8N8sRR:HCM0oRCs:(=RUS;
SNS0LRDC:FRslL0ND
C;S8SSVRD0:FRslsIF82
S;b
SFRs05S
SS7q7)RR:H#MR0D8_FOoH_OPC0RFs58N8s8IH0-ERR84RF0IMF2Rj;S
SSz7maRR:FRk0#_08DHFoOC_POs0FRH5I8R0E-RR48MFI0jFR2S
S2S;
Ns00H0LkChRQQ:aRRs#0H;Mo
0SN0LsHkR0C\N3sMR	\:MRH0CCosR;
RNRR0H0sLCk0Rs\3CPlFCF_M_sINM:\RR0HMCsoC;M
C8MRC0$H0Rv)m_#LNC
;
NEsOHO0C0CksRD#CC_O0)RmvF)VRmLv_NR#CHS#
#0kL$RbCsFFlkH0R#0R#8F_Do_HOP0COFIs5HE80-84RF0IMF2Rj;-
-SlOFbCFMMv0RznXw
S--SsbF0
R5-S-SSRSmRF:Rk#0R0D8_FOoH;-
-SSSSQ:jRRRHM#_08DHFoO-;
-SSSSRQ4:MRHR8#0_oDFH
O;-S-SSRS1RH:RM0R#8F_Do
HO-S-SS
2;-C-SMO8RFFlbM0CM;
S
SMOF#M0N0CREGRR:#H0sMjo5RR0F4R62:"=Rjd4.c(6nUAgqBw7 "
;
SMVkOF0HMFRslL0NDCCsN085NCLDRs:RFNl0L;DCRRI,LD,RC:MRR0HMCsoC2CRs0MksRs#0HRMo=">Rs0FlNCLDs8CN"
;
SMVkOF0HMkRVMNOPDF5L0l0FDCHM_RV,DNFI8_8sVE,RHNoE8_8sVL,RHR0,M0LH#RR:HCM0o2CsR0sCkRsM#H0sMHoR#S
SO#FM00NMRb0FRH:RMo0CC:sR=FRL0l0FDCHM_+VRRHML0-#RR
4;SNSPsLHNDHCR,,R[RRP,L#bFRH:RMo0CC
s;SFSOMN#0M00RFEbON:sRR0HMCsoCRR:=M0LH#RR/cRR-4S;
SsPNHDNLCkRLVRR:#H0sM0o5FEbON8sRF0IMF2Rj;L
SCMoH
HSSVF5L0l0FDCHM_<VRRIDFNs88_FVRsFR0bRR>EEHoNs88_RV20MEC
SSS[=R:R
j;SPSSRR:=jS;
SbSLF:#R=;Rj
SSSVRFsHMRHR0LF0DFlH_MCVFR0Rb0FRFRDFSb
SHSSVRRH<FRDI8N8sR_VFHsRRE>RHNoE8_8sVER0CSM
SSSSH8VRV5D0L2H0R'=R40'RE
CMSSSSSRSP:P=RR.+R*;*[
SSSSMSC8VRH;S
SSDSC#SC
SSSSH0VRNCLD55H2L2H0R'=R40'RE
CMSSSSSRSP:P=RR.+R*;*[
SSSSMSC8VRH;S
SSMSC8VRH;S
SSRS[:[=RR4+R;RRRRR--MLklCFsRVHRL0O#RFCDDO80CRS
SSVSH5=[RRRc20MECRR--CsPC$RRcI8CRkRlbHFM0RONRENNsOs0C
SSSSRS[:j=R;S
SSLSSkLV5b2F#RR:=E5CGP
2;SSSSSFLb#=R:RFLb#RR+4S;
SSSSP=R:R
j;SSSSCRM8H
V;SCSSMD8RF;Fb
SSSskC0sLMRk
V;SDSC#SC
SCSs0MksRlsF0DNLCNsC8N50L,DCR0LF0DFlH_MCVL,RHR0,M0LH#
2;SMSC8VRH;C
SMV8Rk0MOHRFMVOkMP;ND
O
SF0M#NRM0L0F0FHlpM:CRR0HMCsoCRR:=5IDFNs88/24n*;4n
FSOMN#0ML0RFF00lpd.HRMC:MRH0CCos=R:RF5DI8N8s./d2.*d;O
SF0M#NRM0EEHopCHMRH:RMo0CC:sR=ER5HNoE8/8s4*n24
n;SMOF#M0N0HREo.EdpCHMRH:RMo0CC:sR=ER5HNoE8/8sd*.2d
.;SMOF#M0N0HREoFEAss8CRH:RMo0CC:sR=HREoHEpM+CRRR46;O
SF0M#NRM00#sH0CN0_:HRR0HMCsoCRR:=5oEHEsAF8+Cs4F-L0l0FpCHM2n/4RS;
0C$bRL0NRRH#NNss$5R5EEHodH.pM-CRR0LF0dFl.MpHCd2/.R+48MFI0jFR2VRFRlsFFRk0;#
SHNoMDmR1zRa,pamzR0:RN
L;So#HMRND7amz_GNk,mR7zNa_kRG.:0R#8F_Do_HOP0COFIs5HE80-84RF0IMF2Rj;C
Lo
HMRRRRRsVF_bbHCV:RFHsRRRHMjFR0R8IH04E-RMoCC0sNCS
SNs00H0LkC3R\s	NM\VRFRosC#RR:DCNLD#RHR
4;RRRRRRRRNs00H0LkC3R\sFClPMC_FN_IsRM\FsVRCRo#:NRDLRCDH4#R;R
SLHCoMS
SRosC#b:RHLbCkSV
SbSRFRs0l5Nb
RSRRSSSSQRRRR=>7amz_GNk5,H2
RSRRSSSSmRRRR=>7amz5
H2SSSSS;R2
CSRMo8RCsMCNR0CV_FsbCHb;S

H4V_nR#:H5VREEHodH.pM>CRR0LF0dFl.MpHCo2RCsMCN
0CSCSLo
HMSVSH_L4n:VRHRF5L0l0FpCHMRL=RFF00lpd.H2MCRMoCC0sNCS
SSRL:VRFsLRH0HjMRRR0FI0H8ERR-4CRoMNCs0SC
SNSS0H0sLCk0RQQhaVRFRv)m :6RRLDNCHDR#kRVMNOPDF5L0l0FpCHM,FRDI8N8sE,RHNoE8,8sR0LH,.Rd2S;
SCSLo
HMSSSS) mv6RR:)dmv.
X4SSSSSFSbsl0RN5bRRjRqRR=>q)775,j2
SSSSSSSS4SqRR=>q)775,42
SSSSSSSS.SqRR=>q)775,.2
SSSSSSSSdSqRR=>q)775,d2
SSSSSSSScSqRR=>q)775,c2
SSSSSSSSRSmRR=>1amz55j2L2H0
SSSSSSSS;S2
SSSCRM8oCCMsCN0R
L;SMSC8CRoMNCs0HCRVn_4LS;
S_HV4:nLRRHV50LF0pFlHRMC>FRL0l0FdH.pMRC2oCCMsCN0
SSSLV:RFLsRHH0RMRRj0IFRHE80R4-RRMoCC0sNCS
SS0SN0LsHkR0CQahQRRFV) mvcRR:DCNLD#RHRMVkODPN50LF0pFlH,MCRIDFNs88,HREo8EN8Rs,L,H0R24n;S
SSoLCHSM
S)SSmcv R):Rmnv4XS4
SSSSSsbF0NRlbRR5RRqj=q>R757)j
2,SSSSSSSSSRq4=q>R757)4
2,SSSSSSSSSRq.=q>R757).
2,SSSSSSSSSRqd=q>R757)d
2,SSSSSSSSSRmR=1>Rm5zajL25H
02SSSSSSSSS
2;SCSSMo8RCsMCNR0CLS;
S8CMRMoCC0sNCVRH_L4n;C
SMo8RCsMCNR0CH4V_n
#;
VSH_#d.:VRHRH5Eo.EdpCHMRL=RFF00lpd.H2MCRMoCC0sNCS
SH4V_nRO:H5VRL0F0FHlpM=CRR0LF0dFl.MpHCo2RCsMCN
0CSLSS:FRVsHRL0MRHR0jRFHRI8R0E-RR4oCCMsCN0
SSSS_HV4H:RVNR58I8sHE80R4=R2CRoMNCs0SC
SSSSNs00H0LkChRQQFaRVmR)vR 4:NRDLRCDHV#RkPMONLD5FF00lMpHCD,RF8IN8Rs,EEHoNs88,HRL04,Rn
2;SSSSLHCoMS
SS)SSm4v R):Rmnv4XS4
SSSSSFSbsl0RN5bRRjRqRR=>q)775,j2
SSSSSSSSqSS4>R=R''j,S
SSSSSSSSSq=.R>jR''S,
SSSSSSSSSRqd='>Rj
',SSSSSSSSSRSmRR=>1amz55j2L2H0
SSSSSSSS;S2
SSSS8CMRMoCC0sNCVRH_
4;SSSSH.V_:VRHR85N8HsI8R0E=2R.RMoCC0sNCS
SSNSS0H0sLCk0RQQhaVRFRv)m :.RRLDNCHDR#kRVMNOPDF5L0l0FpCHM,FRDI8N8sE,RHNoE8,8sR0LH,nR42S;
SLSSCMoH
SSSSmS)vR .:mR)vX4n4S
SSSSSSsbF0NRlbRR5RRqj=q>R757)j
2,SSSSSSSSS4SqRR=>q)775,42
SSSSSSSSqSS.>R=R''j,S
SSSSSSSSSq=dR>jR''S,
SSSSSSSSSRmR=1>Rm5zajL25H
02SSSSSSSSS
2;SSSSCRM8oCCMsCN0R_HV.S;
SHSSV:_dRRHV58N8s8IH0=ERRRd2oCCMsCN0
SSSS0SN0LsHkR0CQahQRRFV) mvdRR:DCNLD#RHRMVkODPN50LF0pFlH,MCRIDFNs88,HREo8EN8Rs,L,H0R24n;S
SSCSLo
HMSSSSSv)m :dRRv)m44nX
SSSSSSSb0FsRblNRR5Rq=jR>7Rq7j)52S,
SSSSSSSSSRq4=q>R757)4
2,SSSSSSSSS.SqRR=>q)775,.2
SSSSSSSSqSSd>R=R''j,S
SSSSSSSSSm=RR>mR1zja52H5L0S2
SSSSS;S2
SSSS8CMRMoCC0sNCVRH_
d;SSSSHcV_:VRHRE55HNoE8-8sL0F0FHlpM<CRR24nR8NMR85N8HsI8R0E>c=R2o2RCsMCN
0CSSSSS0N0skHL0QCRhRQaF)VRmcv RD:RNDLCRRH#VOkMP5NDL0F0FHlpMRC,DNFI8,8sRoEHE8N8sL,RHR0,4;n2
SSSSoLCHSM
SSSS) mvcRR:)4mvn
X4SSSSSbSSFRs0lRNb5qRRj>R=R7q7)25j,S
SSSSSSSSSq=4R>7Rq74)52S,
SSSSSSSSSRq.=q>R757).
2,SSSSSSSSSdSqRR=>q)775,d2
SSSSSSSSmSSR>R=Rz1ma25j50LH2S
SSSSSS2SS;S
SSMSC8CRoMNCs0HCRV;_c
SSSS_HV6H:RV5R5Ns88I0H8E=R>RR62NRM85oEHE8N8sRR-L0F0FHlpM>CR=nR42o2RCsMCN
0CSSSSS0N0skHL0QCRhRQaF)VRm6v RD:RNDLCRRH#VOkMP5NDL0F0FHlpMRC,DNFI8,8sRoEHE8N8sL,RHR0,d;.2
SSSSoLCHSM
SSSS) mv6RR:)dmv.
X4SSSSSbSSFRs0lRNb5qRRj>R=R7q7)25j,S
SSSSSSSSSq=4R>7Rq74)52S,
SSSSSSSSSRq.=q>R757).
2,SSSSSSSSSdSqRR=>q)775,d2
SSSSSSSSqSSc>R=R7q7)25c,S
SSSSSSSSSm=RR>mR1zja52H5L0S2
SSSSSSSS2S;
SCSSMo8RCsMCNR0CH6V_;S
SS8CMRMoCC0sNC;RL
CSSMo8RCsMCNR0CH4V_n
O;SVSH_84n:VRHRF5L0l0FpCHMRL>RFF00lpd.H2MCRMoCC0sNCS
SS_HVNI8sHE80:VRHR85N8HsI8R0E>2RcRMoCC0sNCS
SS:SLRsVFR0LHRRHMjFR0R8IH0-ERRo4RCsMCN
0CSSSSS_HVcH:RV5R5EEHoNs88-0LF0DFlHRMC<nR42MRN8NR58I8sHE80RR>=cR22oCCMsCN0
SSSSNSS0H0sLCk0RQQhaVRFRv)m :cRRLDNCHDR#kRVMNOPDF5L0l0FpCHM,FRDI8N8sE,RHNoE8,8sR0LH,nR42S;
SSSSLHCoMS
SSSSS) mvcRR:)4mvn
X4SSSSSSSSb0FsRblNRq5Rj>R=R7q7)25j,S
SSSSSSSSSSRq4=q>R757)4
2,SSSSSSSSSqSS.>R=R7q7)25.,S
SSSSSSSSSSRqd=q>R757)d
2,SSSSSSSSSmSSRR=>1amz55j2L2H0
SSSSSSSSSSS2S;
SSSSCRM8oCCMsCN0R_HVcS;
SCSSMo8RCsMCNR0CLS;
SMSC8CRoMNCs0HCRV8_Ns8IH0
E;SHSSV8_N8HsI8:0ERRHV58N8s8IH0<ER=2RcRMoCC0sNCS
SS:SLRsVFR0LHRRHMjFR0R8IH0-ERRo4RCsMCN
0CSSSSS_HV4H:RVNR58I8sHE80R4=R2CRoMNCs0SC
SSSSS0N0skHL0QCRhRQaF)VRm4v RD:RNDLCRRH#VOkMP5NDL0F0FHlpMRC,DNFI8,8sRoEHE8N8sL,RHR0,4;n2
SSSSCSLo
HMSSSSSmS)vR 4:mR)vX4n4S
SSSSSSFSbsl0RN5bRRjRqRR=>q)775,j2
SSSSSSSSSSSq=4R>jR''S,
SSSSSSSSS.SqRR=>',j'
SSSSSSSSSSSq=dR>jR''S,
SSSSSSSSSRSmRR=>1amz55j2L2H0
SSSSSSSS2SS;S
SSCSSMo8RCsMCNR0CH4V_;S
SSHSSV:_.RRHV58N8s8IH0=ERRR.2oCCMsCN0
SSSSNSS0H0sLCk0RQQhaVRFRv)m :.RRLDNCHDR#kRVMNOPDF5L0l0FpCHM,FRDI8N8sE,RHNoE8,8sR0LH,nR42S;
SSSSLHCoMS
SSSSS) mv.RR:)4mvn
X4SSSSSSSSb0FsRblNRR5Rq=jR>7Rq7j)52S,
SSSSSSSSS4SqRR=>q)775,42
SSSSSSSSSSSq=.R>jR''S,
SSSSSSSSSdSqRR=>',j'
SSSSSSSSSSSm=RR>mR1zja52H5L0S2
SSSSSSSSS
2;SSSSS8CMRMoCC0sNCVRH_
.;SSSSS_HVdH:RVNR58I8sHE80Rd=R2CRoMNCs0SC
SSSSS0N0skHL0QCRhRQaF)VRmdv RD:RNDLCRRH#VOkMP5NDL0F0FHlpMRC,DNFI8,8sRoEHE8N8sL,RHR0,4;n2
SSSSCSLo
HMSSSSSmS)vR d:mR)vX4n4S
SSSSSSFSbsl0RN5bRRjRqRR=>q)775,j2
SSSSSSSSSSSq=4R>7Rq74)52S,
SSSSSSSSS.SqRR=>q)775,.2
SSSSSSSSSSSq=dR>jR''S,
SSSSSSSSSRSmRR=>1amz55j2L2H0
SSSSSSSS
2;SSSSS8CMRMoCC0sNCVRH_
d;SSSSS_HVcH:RV5R5EEHoNs88-0LF0DFlHRMC<nR42MRN8NR58I8sHE80RR>=cR22oCCMsCN0
SSSSNSS0H0sLCk0RQQhaVRFRv)m :cRRLDNCHDR#kRVMNOPDF5L0l0FpCHM,FRDI8N8sE,RHNoE8,8sR0LH,nR42S;
SSSSLHCoMS
SSSSS) mvcRR:)4mvn
X4SSSSSSSSb0FsRblNRR5Rq=jR>7Rq7j)52S,
SSSSSSSSS4SqRR=>q)775,42
SSSSSSSSSSSq=.R>7Rq7.)52S,
SSSSSSSSSdSqRR=>q)775,d2
SSSSSSSSSSSm=RR>mR1zja52H5L0S2
SSSSS2SS;S
SSCSSMo8RCsMCNR0CHcV_;S
SSMSC8CRoMNCs0LCR;S
SS8CMRMoCC0sNCVRH_8N8s8IH0
E;SMSC8CRoMNCs0HCRVn_48S;
CRM8oCCMsCN0R_HVd;.#
L
S4V:RFIsRRRHM4FR0RH5Eo.EdpCHMRL-RFF00lpd.H-MCd/.2do.RCsMCN
0CS:SLRsVFR0LHRRHMjFR0R8IH0-ERRo4RCsMCN
0CSNSS0H0sLCk0RQQhaVRFRv)m :6RRLDNCHDR#kRVMNOPD*5IdL.+FF00lpd.H,MCRIDFNs88,HREo8EN8Rs,L,H0R2d.;S
SSo#HMRNDbCHb_k8F0:#RR8#0_oDFH
O;SCSLo
HMS)SSm6v R):Rm.vdXS4
SSSSb0FsRblNRR5Rq=jR>7Rq7j)52S,
SSSSSqSS4>R=R7q7)254,S
SSSSSS.SqRR=>q)775,.2
SSSSSSSSRqd=q>R757)d
2,SSSSSSSSq=cR>7Rq7c)52S,
SSSSSmSSR>R=Rz1ma25I50LH2S
SSSSSS
2;SMSC8CRoMNCs0LCR;C
SMo8RCsMCNR0CL
4;
VSH_F4n:VRHRE55HdoE.MpHCRR=RoEHEMpHCN2RM58REEHodH.pM>CRR0LF0dFl.MpHCR22oCCMsCN0
LSS:FRVsHRL0MRHR0jRFHRI8R0E-RR4oCCMsCN0
SSS#MHoNFDRkC0_M:8RR8#0_oDFH
O;SNSS0H0sLCk0RQQhaVRFRv)m :cRRLDNCHDR#kRVMNOPDH5EoFEAss8C-,46RoEHEsAF8-Cs4R6,EEHoNs88,HRL04,Rn
2;SCSLo
HMS)SSmcv R):Rmnv4XS4
SSSSb0FsRblNRq5Rj=RR>7Rq7j)52S,
SSSSSqSS4>R=R7q7)254,S
SSSSSS.SqRR=>q)775,.2
SSSSSSSSRqd=q>R757)d
2,SSSSSSSSm=RR>mR1z5a5EEHodH.pMLC-FF00lpd.H-MCd/.2d4.+2H5L0S2
SSSSS;S2
CSSMo8RCsMCNR0CLS;
CRM8oCCMsCN0R_HV4;nF
VSH_#4n:VRHRE55HdoE.MpHCRR<RoEHEMpHCN2RM58REEHodH.pM>CRR0LF0dFl.MpHCR22oCCMsCN0
LSS:FRVsHRL0MRHR0jRFHRI8R0E-RR4oCCMsCN0
SSS#MHoNFDRkC0_M:8RR8#0_oDFH
O;SNSS0H0sLCk0RQQhaVRFRv)m :6RRLDNCHDR#kRVMNOPDH5EoFEAss8C-,d4RoEHEsAF8-CsdR4,EEHoNs88,HRL0d,R.
2;SCSLo
HMS)SSm6v R):Rm.vdXS4
SSSSb0FsRblNRR5Rq=jR>7Rq7j)52S,
SSSSSqSS4>R=R7q7)254,S
SSSSSS.SqRR=>q)775,.2
SSSSSSSSRqd=q>R757)d
2,SSSSSSSSq=cR>7Rq7c)52S,
SSSSSmSSR>R=Rz1maE55HdoE.MpHCF-L0l0FdH.pM/C2d5.2L2H0
SSSSSSS2S;
S8CMRMoCC0sNC;RL
MSC8CRoMNCs0HCRVn_4#
;
RRRRHIV_HE80:VRHRs50HN#00HC_R6<R2CRoMNCs0RC
RRRRRHRRVk_F0Rj:H5VREEHodH.pM=CRR0LF0dFl.MpHCo2RCsMCN
0CRRRRRRRRRpRRm5zaj<2R=mR1zja52R;
RRRRRCRRMo8RCsMCNR0CHFV_k;0j
RRRRRRRR_HVF4k0:VRHRH5Eo.EdpCHMRL>RFF00lpd.H2MCRMoCC0sNCR
RRRRRRRRRR_HVOCN#4H:RVLR5FF00lMpHCRR=L0F0F.ldpCHM2CRoMNCs0-C
-#SSHNoMDHR8V:VRR8#0_oDFH
O;SRRRLHCoM-
-RRRRRRRRRRRRRHR8V<VR=jR''ERICqMR7R7)<B=Rm_he1_a7pQmtB _eB)am5+d4L0F0FHlpMRC,Ns88I0H8E
2R-R-RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRCRRDR#C';4'
S--RRRRRFRVsH_I8:0ERsVFRHHRMRRj0IFRHE80-o4RCsMCN
0C-R-SRRRRRRRRl0kGsRCC:zRvX
wn-S-SSsbF0NRlb
R5-S-SSRSRm=RR>mRpzja5225H,-
-SSSSRjRQRR=>1amz55j2H
2,-S-SSRSRQ=4R>mR1z4a5225H,-
-SSSSRRR1RR=>8VHV
S--S;S2
R--RRRRRRRRRRRRR8CMRMoCC0sNCFRVsH_I8;0E
RRRRRRRRRRRRpRRm5zaj<2R=mR1zja52ERICqMR7R7)<B=Rm_he1_a7pQmtB _eB)am5+d4L0F0FHlpMRC,Ns88I0H8E
2RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR#CDCmR1z4a52R;
RRRRRRRRRMRC8CRoMNCs0HCRVN_O#;C4
RRRRRRRRRRRHOV_N.#C:VRHRF5L0l0FpCHMRL>RFF00lpd.H2MCRMoCC0sNC-
-SHS#oDMNRV8HV:jRR8#0_oDFH
O;SRRRRoLCH-M
-RRRRRRRRRRRR8RRHjVVRR<='Rj'IMECR7q7)=R<RhBmea_17m_pt_QBea Bm4)56F+L0l0FpCHM,8RN8HsI820ER-
-RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRCCD#R''4;-
-SRRRRVRRFIs_HE80jV:RFHsRRRHMjFR0R8IH04E-RMoCC0sNC-
-SRRRRRRRRkRlGC0sCRR:vwzXn-
-SbSSFRs0lRNb5-
-SSSSRRRmRR=>pamz55j2H
2,-S-SSRSRQ=jR>mR1zja5225H,-
-SSSSR4RQRR=>1amz5542H
2,-S-SSRSR1=RR>HR8V
Vj-S-SS
2;-R-RRRRRRRRRRRRRCRM8oCCMsCN0RsVF_8IH0;Ej
RRRRRRRRRRRRpRRm5zaj<2R=mR1zja52ERICqMR7R7)<B=Rm_he1_a7pQmtB _eB)am5+46L0F0FHlpMRC,Ns88I0H8E
2RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR#CDCmR1z4a52R;
RRRRRRRRRMRC8CRoMNCs0HCRVN_O#;C.
RRRRRRRR8CMRMoCC0sNCVRH_0Fk4R;
RRRRRNRR:FRVsRRIH4MRRR0F5oEHEpd.HRMC-FRL0l0FdH.pMdC-.d2/.R-4oCCMsCN0
S--So#HMRND8VHV4RR:#_08DHFoOC_POs0F5H5Eo.EdpCHMRL-RFF00lpd.H-MCd/.2d4.-RI8FMR0F4
2;SRRRRoLCH-M
-RRRRRRRRRRRR8RRH4VV5RI2<'=RjI'RERCMq)77RB<Rm_he1_a7pQmtB _eB)am5*d.54I+2F+L0l0FdH.pMRC,Ns88I0H8E-2
-RRRRRRRRRRRRRRRRRRRRRRRRRRRRDRC#'CR4
';-R-SRRRRRsVF_8IH0:E4RsVFRHHRMRRj0IFRHE80-o4RCsMCN
0C-R-SRRRRRRRRl0kGsRCC:zRvX
wn-S-SSsbF0NRlb
R5-S-SSRSRm=RR>mRpzIa5225H,-
-SSSSRjRQRR=>pamz54I-225H,-
-SSSSR4RQRR=>1amz54I+225H,-
-SSSSRRR1RR=>8VHV425I
S--S;S2
R--RRRRRRRRRRRRR8CMRMoCC0sNCFRVsH_I840E;R
RRRRRRRRRRRRRpamz5RI2<p=Rm5zaI2-4RCIEM7Rq7<)RRhBmea_17m_pt_QBea Bmd)5.I*5++42L0F0F.ldpCHM,8RN8HsI820E
RRRRRRRRRRRRRRRRRRRRRRRRRRRRDRC#1CRm5zaI2+4;R
RRRRRRMRC8CRoMNCs0NCR;R
RRRRR
RRRRRRRR_HVD0N#4Rn:H5VR5oEHEpd.HRMC=HREoHEpMRC2NRM85oEHEpd.HRMC-FRL0l0FdH.pM>CRR2nd2CRoMNCs0-C
-#SSHNoMDHR8VRV.:0R#8F_Do;HO
RSRRCRLo
HM-R-RRRRRRRRRRRRR8VHV.=R<R''jRCIEM7Rq7<)RRhBmea_17m_pt_QBea BmE)5HAoEFCs8s6-4,8RN8HsI820ER-
-RRRRRRRRRRRRRRRRRRRRRRRRRRRRR#CDC4R''-;
-RSRRRRRV_FsI0H8ER.:VRFsHMRHR0jRFHRI8-0E4CRoMNCs0-C
-RSRRRRRRlRRksG0C:CRRXvzw-n
-SSSb0FsRblNR-5
-SSSSmRRR>R=RzpmaE55HdoE.MpHCF-L0l0FdH.pMdC-.d2/.H252-,
-SSSSQRRj>R=RzpmaE55HdoE.MpHCF-L0l0FdH.pMdC-.d2/.2-45,H2
S--SRSSRRQ4=1>Rm5za5oEHEpd.H-MCL0F0F.ldpCHM2./d225H,-
-SSSSRRR1RR=>8VHV.-
-S2SS;-
-RRRRRRRRRRRRRMRC8CRoMNCs0VCRFIs_HE80.R;
RRRRRRRRRpRRm5za5oEHEpd.H-MCL0F0F.ldpCHM-2d./2d.RR<=pamz5H5Eo.EdpCHM-0LF0dFl.MpHC.-d2./d-R42
SSSSESICqMR7R7)<mRBh1e_ap7_mBtQ_Be a5m)EEHoA8FsC4s-6N,R8I8sHE802R
RRRRRRRRRRRRRRRRRRDRC#1CRm5za5oEHEpd.H-MCL0F0F.ldpCHM2./d2R;
RRRRRCRRMo8RCsMCNR0CHDV_N4#0n
;
RRRRRRRRHDV_Nd#0.H:RV5R5EEHodH.pM<CRRHREoHEpMRC2NRM85oEHEpd.HRMC-FRL0l0FdH.pM>CRR2nd2CRoMNCs0-C
-#SSHNoMDHR8VRVd:0R#8F_Do;HO
RSRRCRLo
HM-R-RRRRRRRRRRRRR8VHVd=R<R''jRCIEM7Rq7<)RRhBmea_17m_pt_QBea BmE)5HAoEFCs8s4-d,8RN8HsI820ER-
-RRRRRRRRRRRRRRRRRRRRRRRRRRRRR#CDC4R''-;
-RSRRRRRV_FsI0H8ERd:VRFsHMRHR0jRFHRI8-0E4CRoMNCs0-C
-RSRRRRRRlRRksG0C:CRRXvzw-n
-SSSb0FsRblNR-5
-SSSSmRRR>R=RzpmaE55HdoE.MpHCF-L0l0FdH.pMdC-.d2/.H252-,
-SSSSQRRj>R=RzpmaE55HdoE.MpHCF-L0l0FdH.pMdC-.d2/.2-45,H2
S--SRSSRRQ4=1>Rm5za5oEHEpd.H-MCL0F0F.ldpCHM2./d225H,-
-SSSSRRR1RR=>8VHVd-
-S2SS;-
-RRRRRRRRRRRRRMRC8CRoMNCs0VCRFIs_HE80dR;
RRRRRRRRRpRRm5za5oEHEpd.H-MCL0F0F.ldpCHM-2d./2d.RR<=pamz5H5Eo.EdpCHM-0LF0dFl.MpHC.-d2./d-R42
SSSSESICqMR7R7)<mRBh1e_ap7_mBtQ_Be a5m)EEHoA8FsCds-4N,R8I8sHE802R
RRRRRRRRRRRRRRRRRRDRC#1CRm5za5oEHEpd.H-MCL0F0F.ldpCHM2./d2R;
RRRRRCRRMo8RCsMCNR0CHDV_Nd#0.
;
RRRRRRRRHFV_k:0.RRHV5oEHEsAF8RCs-FRL0l0FpCHMRn<Rco2RCsMCN
0CRRRRRRRRRRRRRmR7zNa_k<GR=VR8DI0RERCM5RRRR75q7>)RRhBmea_17m_pt_QBea BmE)5HAoEFCs8sN,R8I8sHE802R2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRF5sRq)77RB<Rm_he1_a7pQmtB _eB)am50LF0pFlH,MCR8N8s8IH02E22R
RRRRRRRRRRRRRRRRRRRRRRRRRR#CDCmRpzja52R;
RRRRRCRRMo8RCsMCNR0CHFV_k;0.
RRRRRRRR_HVFdk0:VRHRH5EoFEAss8CRL-RFF00lMpHCRR>nRd2oCCMsCN0
RRRRRRRRRRRR7RRm_zaNRkG<8=RVRD0IMECRR5RRqR57R7)>mRBh1e_ap7_mBtQ_Be a5m)EEHoA8FsCRs,Ns88I0H8E
22RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRsRFR75q7<)RRhBmea_17m_pt_QBea BmL)5FF00lMpHCN,R8I8sHE802
22RRRRRRRRRRRRRRRRRRRRRRRRRCRRDR#Cpamz5H5Eo.EdpCHM-0LF0dFl.MpHC.-d2./d2R;
RRRRRCRRMo8RCsMCNR0CHFV_k;0d
RRRRMRC8CRoMNCs0HCRVH_I8;0E
RRR
RRRRVRH_8IH0:EjRRHV5H0s#00NCR_H>6=R2CRoMNCs0RC
RRRRRHRRVN_O#:C4RRHV50LF0pFlHRMC=FRL0l0FdH.pMRC2oCCMsCN0
RRRRRRRRRRR7amz_GNkRR<=1amz5Rj2IMECRR5RRqR57R7)<B=Rm_he1_a7pQmtB _eB)am5+d4L0F0FHlpMRC,Ns88I0H8ER22
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRMRN8qR57R7)>B=Rm_he1_a7pQmtB _eB)am50LF0pFlH,MCR8N8s8IH02E22R
RRRRRRRRRRRRRRRRRRRRRRRRRR#CDCFRsl0Fk'05FE#CsRR=>'2Z';R
RRRRRRMRC8CRoMNCs0HCRVN_O#;C4
RRRRRRRR_HVOCN#.H:RVLR5FF00lMpHCRR>L0F0F.ldpCHM2CRoMNCs0RC
RRRRRRRRRmR7zNa_k<GR=mR1zja52ERIC5MRRRRR57q7)=R<RhBmea_17m_pt_QBea Bm4)56F+L0l0FpCHM,8RN8HsI820E2RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRSMRN8qR57R7)>B=Rm_he1_a7pQmtB _eB)am50LF0pFlH,MCR8N8s8IH02E22R
RRRRRRRRRRRRRRRRRRRRRRRRRR#CDCFRsl0Fk'05FE#CsRR=>'2Z';R
RRRRRRMRC8CRoMNCs0HCRVN_O#;C.
RRRRRRRR:NjRsVFRHIRMRR405FREEHodH.pMLC-FF00lpd.H-MCd/.2do.RCsMCN
0CRRRRRRRRRRRRRmR7zNa_k<GR=mR1zIa52ERIC5MRRRRR57q7)=R<RhBmea_17m_pt_QBea Bmd)5.I*5++42R0LF0dFl.MpHC,-4R8N8s8IH02E2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR8NMR75q7>)R=mRBh1e_ap7_mBtQ_Be a5m)dI.*+0LF0dFl.MpHCN,R8I8sHE802
22RRRRRRRRRRRRRRRRRRRRRRRRRRRRRDRC#sCRFklF0F'50sEC#>R=R''Z2R;
RRRRRCRRMo8RCsMCNR0CN
j;RRRRRRRRH#V_k.bd:VRHRE55HdoE.MpHCRR=RoEHEMpHCN2RM58REEHodH.pM-CRR0LF0dFl.MpHCRR>n2d2RMoCC0sNCR
RRRRRRRRRRRRR7amz_GNkRR<=1amz5H5Eo.EdpCHM-0LF0dFl.MpHCd2/.
2RSRSSRSSSSCIEMRR5R5RRq)77RR<=Bemh_71a_tpmQeB_ mBa)H5EoFEAss8C,8RN8HsI820E2R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRNRM857q7)=R>RhBmea_17m_pt_QBea BmE)5HAoEFCs8s6-4,8RN8HsI820E2R2
RRRRRRRRRRRRRRRRRRRRRRRRRCRRDR#CsFFlk50'FC0Es=#R>ZR''
2;RRRRRRRRCRM8oCCMsCN0R_HV#dkb.R;
RRRRRHRRVk_#b:4nRRHV5H5Eo.EdpCHMRR<REEHopCHM2MRN8ER5HdoE.MpHCRR-L0F0F.ldpCHMRn>RdR22oCCMsCN0
RRRRRRRRRRRR7RRm_zaNRkG<1=Rm5za5oEHEpd.H-MCL0F0F.ldpCHM2./d2SR
SRSRSSSSIMECRR5RRqR57R7)<B=Rm_he1_a7pQmtB _eB)am5oEHEsAF8,CsR8N8s8IH02E2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRNRRM58Rq)77RR>=Bemh_71a_tpmQeB_ mBa)H5EoFEAss8C-,d4R8N8s8IH02E22R
RRRRRRRRRRRRRRRRRRRRRRRRRRDRC#sCRFklF0F'50sEC#>R=R''Z2R;
RRRRRCRRMo8RCsMCNR0CH#V_knb4;R
RRRRRRVRH_IDF:VRHRF5L0l0FpCHMRj>R2CRoMNCs0RC
RRRRRRRRRmR7zNa_k<GR=VR8DI0RERCM5RRR57q7)RR<Bemh_71a_tpmQeB_ mBa)F5L0l0FpCHM,8RN8HsI820E2R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRSFRRsqR57R7)>mRBh1e_ap7_mBtQ_Be a5m)EEHoA8FsCRs,Ns88I0H8E222
RRRRRRRRRRRRRRRRRRRRRRRR#CDCFRsl0Fk'05FE#CsRR=>'2Z';R
RRRRRRMRC8CRoMNCs0HCRVF_DIR;
RRRRRHRRVF_DIRj:H5VRL0F0FHlpM<CRRR42oCCMsCN0
RRRRRRRRRRR7amz_GNkRR<=80VDRCIEMqR57R7)>mRBh1e_ap7_mBtQ_Be a5m)EEHoA8FsCRs,Ns88I0H8E
22RRRRRRRRRRRRRRRRRRRRRRRRCCD#RlsFF'k05EF0CRs#='>RZ;'2
RRRRRRRR8CMRMoCC0sNCVRH_IDFjR;
RRRRCRM8oCCMsCN0R_HVI0H8E
j;
8CMRONsECH0Os0kCCR#D0CO_v)m;D

HNLssH$RC;CC
Ck#RCHCC03#8F_Do_HO4c4n3DND;#
kCCRHC#C30D8_FOoH_HNs0NE3D
D;kR#CHCCC38#0_oDFHkO_Mo#HM3C8N;DD
Ck#RsIF	C3oMObN	CNo3DND;D

HNLssk$RMHH#lk;
#kCRMHH#lO3PFFlbM0CM#D3ND
;
CHM00)$RmHvR#o
SCsMCH5OR
SSSVHNlD:$RRs#0HRMo:"=RN"M$;S
SS8IH0:ERR0HMCsoCRR:=cS;
S8SN8HsI8R0E:MRH0CCos=R:R
(;SDSSF8IN8:sRR0HMCsoCRR:=jS;
SHSEo8EN8:sRR0HMCsoCRR:=(
U;S0SSNCLDRs:RFNl0L;DC
SSS80VDRs:RFFlIsS8
2S;
b0FsRS5
S7Sq7:)RRRHM#_08DHFoOC_POs0FR85N8HsI8R0E-RR48MFI0jFR2S;
SmS7z:aRR0FkR8#0_oDFHPO_CFO0sIR5HE80R4-RRI8FMR0FjS2
S
2;
0SN0LsHkR0C\N3sMR	\:MRH0CCosR;
RNRR0H0sLCk0Rs\3CPlFCF_M_sINM:\RR0HMCsoC;M
C8MRC0$H0Rv)m;N

sHOE00COkRsC#CCDO)0_mFvRVmR)v#RH
FSOlMbFCRM0)_mvLCN#
oSSCsMCH5OR
SSSS8IH0:ERR0HMCsoC;S
SS8SN8HsI8R0E:MRH0CCosS;
SDSSF8IN8:sRR0HMCsoC;S
SSHSEo8EN8:sRR0HMCsoC;S
SSNS0LRDC:FRslL0ND
C;SSSS80VDRs:RFFlIsS8
S
2;SFSbs50R
SSSS7q7)RR:H#MR0D8_FOoH_OPC0RFs58N8s8IH0-ERR84RF0IMF2Rj;S
SSmS7z:aRR0FkR8#0_oDFHPO_CFO0sIR5HE80R4-RRI8FMR0FjS2
S;S2
MSC8FROlMbFC;M0
O
SF0M#NRM0MR0L:MRH0CCos=R:R;4n
V
Sk0MOHRFM#s0N0l)FpCHMR0sCkRsMHCM0oRCsHS#
SsPNHDNLCHR#x:CRR0HMCsoC;S
SO#FM00NMRFLDOH	#x:CRR0HMCsoCRR:=MR0L*cRn;L
SCMoH
HSSVDR5F8IN8lsRFL8RD	FO#CHx2RR=R0jRE
CMSsSSCs0kMFRDI8N8sRR+LODF	x#HCS;
S#CDCS
SS0sCkRsM5F5DI8N8sRR+LODF	x#HCRR-4/2RRFLDOH	#xRC2*DRLF#O	H;xC
CSSMH8RVS;
CRM8VOkM0MHFRN#0sF0)lMpHC
;
SMOF#M0N0DRLF#O	HRxC:MRH0CCos=R:RRnc*0RMLS;
O#FM00NMRlDHqs88RH:RMo0CC:sR=0R#N)s0FHlpMRC;
FSOMN#0MM0RLF_sls_VN:ORR0HMCsoCRR:=5oEHE8N8sRR-DqHl8R8s+2R4/DRLF#O	H;xC
FSOMN#0MD0RC_V0s_FlVOsNRH:RMo0CC:sR=ER5HNoE8R8s-HRDl8q8sRR+4l2RFL8RD	FO#CHx;S

0C$bRL0ND8C_FRk0HN#Rs$sNRL5M_lsF_NVsOR+48MFI0jFR2VRFRlsFI8Fs;S

#MHoN8DRF_k0sRFl:NR0L_DC80Fk;C
Lo
HM
VSH_oLH):mvRRHV5oEHE8N8sRR-DNFI8R8s+RR4>DRLF#O	H2xCRMoCC0sNCS
S#MHoN8DRF_k0V#Hs07,Rm_zaNRkG:FRslsIF8S;
So#HMRNDq)77_GNk,7Rq7V)_R#:R0D8_FOoH_OPC0RFs58N8s8IH0-ERR84RF0IMF2Rj;L
SCMoH
S
SV_FsbCHb:FRVsRRHHjMRRR0FNs88I0H8ER-4oCCMsCN0
SSSNs00H0LkC3R\s	NM\VRFRosC#:qRRLDNCHDR#;Rj
SSSNs00H0LkC3R\s	NM\VRFRosC#:ARRLDNCHDR#;R4
RRRRRRRRRRRR0N0skHL0\CR3lsCF_PCMIF_N\sMRRFVs#CoqRR:DCNLD#RHR
4;RRRRRRRRRRRRNs00H0LkC3R\sFClPMC_FN_IsRM\FsVRCAo#RD:RNDLCRRH#4S;
SoLCHSM
SCSso:#qRbbHCVLk
SSSb0FsRblN5S
SSRSSQ>R=R7q7)25H,S
SSSSRR=mR>7Rq7V)_5
H2SSSSS
2;
SSSs#CoAb:RHLbCkSV
SFSbsl0RN
b5SSSSSRRQ=q>R7_7)V25H,S
SSSSRR=mR>7Rq7N)_kHG52S
SS2SS;S
SCRM8oCCMsCN0RsVF_bbHC
;
SmS)v( 4R):RmLv_N
#CSoSSCsMCHlORN
b5SSSSI0H8ESRS=I>RHE80,S
SS8SN8HsI8R0ER>S=R8N8s8IH0RE,
SSSSIDFNs88RSRR=D>RF8IN8
s,SSSSEEHoNs88RSRR=D>RH8lq84s-,S
SSNS0LRDCR=RS>NR0L,DC
SSSSD8V0RRRS>S=RD8V0S
SSS2
SFSbsl0RN5bRR7Rq7=)R>7Rq7V)_,SR
SSSSSz7ma>R=Rk8F0H_Vs
#0SSSSSS2;
S
S80Fk_lsF5Rj2<8=RF_k0V#Hs0ERIC5MRq)77_GNkRR>=Bemh_71a_tpmQeB_ mBa)F5DI8N8sN,R8I8sHE802S2
SSSSSRSSRDRC#8CRV;D0
S
SV_FsDbFF:FRVsRRHH4MRRR0FMsL_FVl_sRNOoCCMsCN0
SSS#MHoN8DRF_k0#o0NCRR:sIFlF;s8
LSSCMoH
SSS) mv6RR:)_mvLCN#
SSSoCCMsRHOl5Nb
SSSS8IH0SERSR=>I0H8ES,
SNSS8I8sHE80R=RS>8RN8HsI8,0ERS
SSFSDI8N8sRRRSR=>DqHl8R8s+HR5-*42LODF	x#HCS,
SESSHNoE8R8sR=RS>HRDl8q8sRR+HD*LF#O	H-xC4
,RSSSS0DNLCRRRSR=>0DNLCS,
S8SSVRD0RSRS=8>RV
D0S2SS
SSSb0FsRblNRR5Rq)77RR=>q)77_RV,
SSSS7SSmRza=8>RF_k0#o0NCS
SS2SS;
S
S8SSF_k0s5FlH<2R=FR8k#0_0CNoRCIEMqR57_7)NRkG>B=Rm_he1_a7pQmtB _eB)am5lDHqs88+-5H4L2*D	FO#CHx,8RN8HsI820E2S
SSSSSSRSRR#CDCFR8ks0_FHl5-;42
CSSMo8RCsMCNR0CV_FsDbFF;

SSVSH_x#HCH:RVDR5C_V0s_FlVOsNRj>R2CRoMNCs0SC
SHS#oDMNRk8F00_#NRoC:FRslsIF8S;
SoLCHSM
SmS)vR 6:mR)vN_L#SC
SCSoMHCsONRlbS5
SISSHE80R=SS>HRI8,0E
SSSS8N8s8IH0RERSR=>Ns88I0H8E
,RSSSSDNFI8R8sR=RS>HRDl8q8sRR+MsL_FVl_s*NOLODF	x#HCS,
SESSHNoE8R8sR=RS>HREo8EN8Rs,
SSSSL0NDRCRR>S=RL0ND
C,SSSS80VDRSRRSR=>80VD
SSS2S
SSsbF0NRlbRR5R7q7)>R=R7q7),_VRS
SSSSS7amzRR=>80Fk_N#0oSC
SSSS2
;SSS
SSk8F0F_slL5M_lsF_NVsO2+4RR<=80Fk_lsF5_MLs_FlVOsN2S
SSSSSSSSSSCIEMqR57_7)NRkG<mRBh1e_ap7_mBtQ_Be a5m)DqHl8+8sMsL_FVl_s*NOLODF	x#HCN,R8I8sHE802S2
SSSSSRSSRSRSRRRRCCD#Rk8F00_#N;oC
SS
SmS7zNa_k<GR=VR8DI0RERCM57q7)k_NGRR>Bemh_71a_tpmQeB_ mBa)H5Eo8EN8Rs,Ns88I0H8E
22SSSSSRSSCCD#Rk8F0F_slL5M_lsF_NVsO2+4;S
SCRM8oCCMsCN0R_HV#CHx;

SSVSH_HM#xRC:H5VRD0CV_lsF_NVsORR=jo2RCsMCN
0CS7SSm_zaNRkG<8=RVRD0IMECR75q7N)_k>GRRhBmea_17m_pt_QBea BmE)5HNoE8,8sR8N8s8IH02E2
SSSSSSSR#CDCFR8ks0_FMl5LF_sls_VN;O2
CSSMo8RCsMCNR0CHMV_#CHx;S

SsVF_bbHCV:RFHsRRRHMjFR0R8IH04E-RMoCC0sNCS
SS0N0skHL0\CR3MsN	F\RVCRso:#RRLDNCHDR#;R.
RRRRRRRRRRRR0N0skHL0\CR3lsCF_PCMIF_N\sMRRFVs#CoRD:RNDLCRRH#4S;
SCRLo
HMSRSSs#Co:HRbbkCLVS
SSbSRFRs0l5Nb
RSSRSRSSRSRQ>R=Rz7mak_NG25H,S
SRSRRSRSSR=mR>mR7zHa52S
SSSSSR
2;SCSRMo8RCsMCNR0CV_FsbCHb;S

CRM8oCCMsCN0R_HVL)Hom
v;
VSH_N#lDmD)vH:RVER5HNoE8R8s-FRDI8N8sRR+4=R<RFLDOH	#xRC2oCCMsCN0
#SSHNoMD7Rq7V)_R#:R0D8_FOoH_OPC0RFs58N8s8IH0-ERR84RF0IMF2Rj;L
SCMoH
VSSFbs_H:bCRsVFRHHRMRRj0NFR8I8sHE80-o4RCsMCN
0CS0SN0LsHkR0C\N3sMR	\FsVRCqo#RD:RNDLCRRH#jS;
S0N0skHL0\CR3lsCF_PCMIF_N\sMRRFVs#CoqRR:DCNLD#RHR
4;SCSLo
HMSsSSCqo#:HRbbkCLVS
SSFSbsl0RN
b5SSSSS=QR>7Rq7H)52S,
SSSSm>R=R7q7)5_VHS2
S2SS;S
SCRM8oCCMsCN0RsVF_bbHC
;
Sv)m :6RRv)m_#LNCS
SSCSoMHCsONRlbS5
SSSSSHSI8R0ES>S=R8IH0
E,RSRSSSSSS8N8s8IH0RERRR=>Ns88I0H8E
,RSSSSSDSSF8IN8RsRR>S=RIDFNs88,S
SSSSSSoEHE8N8sRRRSR=>EEHoNs88,S
SSSSSSL0NDRCRR>S=RL0ND
C,SSSSS8SSVRD0RSRS=8>RV
D0SSSSS2SS
SSSSsbF0NRlbRR5R7q7)>R=R7q7),_VRS
SSSSSSz7ma>R=Rz7maS
SSSSS2
;S
MSC8CRoMNCs0HCRVl_#N)DDm
v;
8CMRONsECH0Os0kCCR#D0CO_v)m;



