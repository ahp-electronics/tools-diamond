library verilog;
use verilog.vl_types.all;
entity config_sspi_dat_cnt is
    port(
        por             : in     vl_logic;
        clk             : in     vl_logic;
        sispi           : in     vl_logic;
        csspi           : in     vl_logic;
        sso             : in     vl_logic;
        rst_exe_r       : in     vl_logic;
        cmd_dec_r       : in     vl_logic;
        cmd_inf_r       : in     vl_logic;
        dat_shf_r       : in     vl_logic;
        cmd_dec         : in     vl_logic;
        dat_shf         : in     vl_logic;
        selasr          : in     vl_logic;
        seldsr          : in     vl_logic;
        prog_inst       : in     vl_logic;
        vfy_inst        : in     vl_logic;
        progstatus_ee_o : in     vl_logic;
        readstatus_ee_o : in     vl_logic;
        flash_status    : in     vl_logic;
        sram_read       : in     vl_logic;
        flash_read      : in     vl_logic;
        vfy_reg32_inst  : in     vl_logic;
        inc_inst        : in     vl_logic;
        sf_secty        : in     vl_logic;
        e2_secty        : in     vl_logic;
        read_tag_o      : in     vl_logic;
        protect_shift_o : in     vl_logic;
        jtag_active     : in     vl_logic;
        instruction     : out    vl_logic_vector(7 downto 0);
        sspi_asrce      : out    vl_logic;
        sspi_dsrce      : out    vl_logic;
        sspi_prechg     : out    vl_logic;
        sspi_read_en    : out    vl_logic;
        sspi_wl_read_str: out    vl_logic;
        sspi_wl_read_str_emb: out    vl_logic;
        sspi_vfy_cap    : out    vl_logic;
        sspi_capdr      : out    vl_logic;
        sospi           : out    vl_logic;
        sospi_en        : out    vl_logic;
        ssi_en          : out    vl_logic;
        sso_en          : out    vl_logic;
        sspi_data       : out    vl_logic;
        sspi_addr       : out    vl_logic;
        byte_cnt        : out    vl_logic_vector(1 downto 0);
        byte_bndy       : out    vl_logic;
        sspi_dsr_preload: out    vl_logic;
        sso_active      : out    vl_logic
    );
end config_sspi_dat_cnt;
