library verilog;
use verilog.vl_types.all;
entity TCK_TREE is
    port(
        A               : in     vl_logic;
        Z               : out    vl_logic
    );
end TCK_TREE;
