library verilog;
use verilog.vl_types.all;
entity MPC_CLK_TREE is
    port(
        A               : in     vl_logic;
        Z               : out    vl_logic
    );
end MPC_CLK_TREE;
