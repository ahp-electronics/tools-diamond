-- $Header: //synplicity/map202003lat/mappers/lattice/lib/gen_lava1/dec.vhd#1 $
@ER--7
 B
LDHs$NsR Q  k;
#QCR 3  #_08DHFoO4_4nNc3D
D;
M
C0$H0RB7 R
H#
MoCCOsH5:MRR0HMCsoC:2=U;b

F5s0
R
q:MRHR8#0_oDFHPO_CFO0s-5M4FR8IFM0R;j2
R
1:kRF00R#8F_Do_HOP0COFMs5-84RF0IMF2Rj
;
2
M
C8 R7B
;
NEsOHO0C0CksR_pe7R BF7VR HBR#O

FFlbM0CMRBeB
RRRb0Fs5R
RRRRRXRRRRRRRRRRRRRRRRRRRRRRRRRRRR:RRRkRF0RRR1_a7pQmtB=R:R''42C;
MO8RFFlbM0CM;O

FFlbM0CMR7th
RRRb0Fs5R
RRRRRXRRRRRRRRRRRRRRRRRRRRRRRRRRRR:RRRkRF0RRR1_a7pQmtB=R:R''j2C;
MO8RFFlbM0CM;O

FFlbM0CMRzBB_A1z
RRRb0Fs5R
RRRRRqRjRRRRRRRRRRRRRRRRRRRRRRRRRR:RRRMRHRRRR1_a7pQmtBR;
RRRRRRAjRRRRRRRRRRRRRRRRRRRRRRRRRRRR:HRRMRRRR71a_tpmQ
B;RRRRRQRBhRRRRRRRRRRRRRRRRRRRRRRRRRRRRR:RHRMRRaR17m_pt;QB
RRRR1RRjRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR:R0FkR1RRap7_mBtQ;R
RRRRRBamzRRRRRRRRRRRRRRRRRRRRRRRRR:RRRkRF0RRR1_a7pQmtB
2;CRM8ObFlFMMC0
;

o#HMRNDOsNs$RRR:0R#8F_Do_HOP0COFRs5MR-48MFI0jFRR
2;#MHoNODRF0M#_:4RR8#0_oDFH
O;#MHoNODRF0M#_:jRR8#0_oDFH
O;
oLCHRM
RRRRRzRR4e:RBuBRmR)av5quR>X=RMOF#40_2R;
RRRRRzRR.t:Rhu7RmR)avRqu5=XR>FROM_#0j
2;RRRRRRRRzRd:B_Bz1RzAuam)Ruvq55RqjR2,O#FM0,_4RMOF#40_,5R1jR2,OsNs$25j2R;
RRRRRzRRcV:RFHsRRRHM4FR0R4M-RMoCC0sNCR
RRRRRRRRRRRRRR.Rz_Rp4:BRBzz_1AmRu)vaRqRu5q25H,FROM_#0jO,RN$ss54H-21,R5,H2RsONsH$52
2;RRRRRRRRCRM8oCCMsCN0;C

Mp8Re _7B
;

