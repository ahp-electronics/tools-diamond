library verilog;
use verilog.vl_types.all;
entity LN0_UDP is
    -- This module cannot be connected to from
    -- VHDL because it has unnamed ports.
end LN0_UDP;
