library verilog;
use verilog.vl_types.all;
entity invx16v1mce is
    port(
        A               : in     vl_logic;
        Z               : out    vl_logic
    );
end invx16v1mce;
