library verilog;
use verilog.vl_types.all;
entity US_DEL is
    port(
        A               : in     vl_logic;
        Y               : out    vl_logic
    );
end US_DEL;
