library verilog;
use verilog.vl_types.all;
entity char_test_logic is
    port(
        cout            : out    vl_logic_vector(19 downto 0);
        char_test_mode  : out    vl_logic;
        char_td         : out    vl_logic_vector(9 downto 0);
        testclk_mst     : in     vl_logic;
        testclk         : out    vl_logic;
        bist_rstn       : out    vl_logic;
        do_bist         : out    vl_logic;
        cptdr           : out    vl_logic;
        shdr            : out    vl_logic;
        bistrtcntdone   : out    vl_logic;
        cin             : in     vl_logic_vector(10 downto 0);
        char_mode       : in     vl_logic;
        rd0             : in     vl_logic_vector(9 downto 0);
        rck0            : in     vl_logic;
        tck0            : in     vl_logic;
        ebrd_clk0       : in     vl_logic;
        fb_clk0         : in     vl_logic;
        rlol0           : in     vl_logic;
        rlos_hi0        : in     vl_logic;
        rlos_lo0        : in     vl_logic;
        pci_connect0    : in     vl_logic;
        pci_det_done0   : in     vl_logic;
        rd1             : in     vl_logic_vector(9 downto 0);
        rck1            : in     vl_logic;
        tck1            : in     vl_logic;
        ebrd_clk1       : in     vl_logic;
        fb_clk1         : in     vl_logic;
        rlol1           : in     vl_logic;
        rlos_hi1        : in     vl_logic;
        rlos_lo1        : in     vl_logic;
        pci_connect1    : in     vl_logic;
        pci_det_done1   : in     vl_logic;
        rd2             : in     vl_logic_vector(9 downto 0);
        rck2            : in     vl_logic;
        tck2            : in     vl_logic;
        ebrd_clk2       : in     vl_logic;
        fb_clk2         : in     vl_logic;
        rlol2           : in     vl_logic;
        rlos_hi2        : in     vl_logic;
        rlos_lo2        : in     vl_logic;
        pci_connect2    : in     vl_logic;
        pci_det_done2   : in     vl_logic;
        rd3             : in     vl_logic_vector(9 downto 0);
        rck3            : in     vl_logic;
        tck3            : in     vl_logic;
        ebrd_clk3       : in     vl_logic;
        fb_clk3         : in     vl_logic;
        rlol3           : in     vl_logic;
        rlos_hi3        : in     vl_logic;
        rlos_lo3        : in     vl_logic;
        pci_connect3    : in     vl_logic;
        pci_det_done3   : in     vl_logic;
        plol            : in     vl_logic;
        rx_ch           : in     vl_logic_vector(3 downto 0);
        bist_rssigso    : in     vl_logic;
        ubs_bistcomplete: in     vl_logic;
        bist_flag_local : in     vl_logic_vector(11 downto 0)
    );
end char_test_logic;
