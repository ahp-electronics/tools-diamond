library verilog;
use verilog.vl_types.all;
entity pcs_quad_top is
    port(
        HDINP0          : in     vl_logic;
        HDINN0          : in     vl_logic;
        HDINP1          : in     vl_logic;
        HDINN1          : in     vl_logic;
        HDINP2          : in     vl_logic;
        HDINN2          : in     vl_logic;
        HDINP3          : in     vl_logic;
        HDINN3          : in     vl_logic;
        HDOUTP0         : out    vl_logic;
        HDOUTN0         : out    vl_logic;
        HDOUTP1         : out    vl_logic;
        HDOUTN1         : out    vl_logic;
        HDOUTP2         : out    vl_logic;
        HDOUTN2         : out    vl_logic;
        HDOUTP3         : out    vl_logic;
        HDOUTN3         : out    vl_logic;
        REFCLKP         : in     vl_logic;
        REFCLKN         : in     vl_logic;
        RXREFCLKP       : in     vl_logic;
        RXREFCLKN       : in     vl_logic;
        RESP            : inout  vl_logic;
        VDDIB0          : in     vl_logic;
        VDDIB1          : in     vl_logic;
        VDDIB2          : in     vl_logic;
        VDDIB3          : in     vl_logic;
        VDDOB0          : in     vl_logic;
        VDDOB1          : in     vl_logic;
        VDDOB2          : in     vl_logic;
        VDDOB3          : in     vl_logic;
        VDDAX25         : in     vl_logic;
        VDDRX0          : in     vl_logic;
        VDDRX1          : in     vl_logic;
        VDDRX2          : in     vl_logic;
        VDDRX3          : in     vl_logic;
        VDDTX0          : in     vl_logic;
        VDDTX1          : in     vl_logic;
        VDDTX2          : in     vl_logic;
        VDDTX3          : in     vl_logic;
        VSSRX           : in     vl_logic;
        VSSTX           : in     vl_logic;
        VDDP            : in     vl_logic;
        VSSP            : in     vl_logic;
        iref50_ext_0    : inout  vl_logic;
        iref50_ext_1    : inout  vl_logic;
        iref50_ext_2    : inout  vl_logic;
        iref50_ext_3    : inout  vl_logic;
        iref50_int_0    : inout  vl_logic;
        iref50_int_1    : inout  vl_logic;
        iref50_int_2    : inout  vl_logic;
        iref50_int_3    : inout  vl_logic;
        iref50_ext_in   : inout  vl_logic;
        iref50_int_in   : inout  vl_logic;
        resp_use        : in     vl_logic;
        logic_hi        : out    vl_logic;
        logic_low       : out    vl_logic;
        scb_rate_sel0   : in     vl_logic_vector(1 downto 0);
        scb_rate_sel1   : in     vl_logic_vector(1 downto 0);
        scb_rate_sel2   : in     vl_logic_vector(1 downto 0);
        scb_rate_sel3   : in     vl_logic_vector(1 downto 0);
        scb_tx_ctl_b    : in     vl_logic_vector(7 downto 0);
        scb_tx_ctl_c    : in     vl_logic_vector(7 downto 0);
        scb_tx_ctl_d    : in     vl_logic_vector(7 downto 0);
        scb_rx_ctl_b    : in     vl_logic_vector(7 downto 0);
        scb_rx_ctl_c    : in     vl_logic_vector(7 downto 0);
        scb_rx_ctl_d    : in     vl_logic_vector(7 downto 0);
        scb_rx_ctl_e    : in     vl_logic_vector(7 downto 0);
        scb_rx_ctl_f    : in     vl_logic_vector(7 downto 0);
        scb_rx_ctl_g    : in     vl_logic_vector(7 downto 0);
        scb_rx_ctl_h    : in     vl_logic_vector(7 downto 0);
        scb_cdr_ctl_a0  : in     vl_logic_vector(7 downto 0);
        scb_cdr_ctl_b0  : in     vl_logic_vector(7 downto 0);
        scb_cdr_ctl_c0  : in     vl_logic_vector(7 downto 0);
        scb_cdr_ctl_d0  : in     vl_logic_vector(7 downto 0);
        scb_cdr_ctl_e0  : in     vl_logic_vector(7 downto 0);
        scb_cdr_ctl_f0  : in     vl_logic_vector(7 downto 0);
        scb_cdr_ctl_g0  : in     vl_logic_vector(7 downto 0);
        scb_cdr_ctl_a1  : in     vl_logic_vector(7 downto 0);
        scb_cdr_ctl_b1  : in     vl_logic_vector(7 downto 0);
        scb_cdr_ctl_c1  : in     vl_logic_vector(7 downto 0);
        scb_cdr_ctl_d1  : in     vl_logic_vector(7 downto 0);
        scb_cdr_ctl_e1  : in     vl_logic_vector(7 downto 0);
        scb_cdr_ctl_f1  : in     vl_logic_vector(7 downto 0);
        scb_cdr_ctl_g1  : in     vl_logic_vector(7 downto 0);
        scb_cdr_ctl_a2  : in     vl_logic_vector(7 downto 0);
        scb_cdr_ctl_b2  : in     vl_logic_vector(7 downto 0);
        scb_cdr_ctl_c2  : in     vl_logic_vector(7 downto 0);
        scb_cdr_ctl_d2  : in     vl_logic_vector(7 downto 0);
        scb_cdr_ctl_e2  : in     vl_logic_vector(7 downto 0);
        scb_cdr_ctl_f2  : in     vl_logic_vector(7 downto 0);
        scb_cdr_ctl_g2  : in     vl_logic_vector(7 downto 0);
        scb_cdr_ctl_a3  : in     vl_logic_vector(7 downto 0);
        scb_cdr_ctl_b3  : in     vl_logic_vector(7 downto 0);
        scb_cdr_ctl_c3  : in     vl_logic_vector(7 downto 0);
        scb_cdr_ctl_d3  : in     vl_logic_vector(7 downto 0);
        scb_cdr_ctl_e3  : in     vl_logic_vector(7 downto 0);
        scb_cdr_ctl_f3  : in     vl_logic_vector(7 downto 0);
        scb_cdr_ctl_g3  : in     vl_logic_vector(7 downto 0);
        scb_pll_ctl_a   : in     vl_logic_vector(7 downto 0);
        scb_pll_ctl_b   : in     vl_logic_vector(7 downto 0);
        scb_pll_ctl_c   : in     vl_logic_vector(7 downto 0);
        scb_pll_ctl_d   : in     vl_logic_vector(7 downto 0);
        scb_pll_ctl_e   : in     vl_logic_vector(7 downto 0);
        scb_pll_ctl_f   : in     vl_logic_vector(7 downto 0);
        scb_pll_ctl_g   : in     vl_logic_vector(7 downto 0);
        scb_ibias_a     : in     vl_logic_vector(7 downto 0);
        scb_bstsds_a    : in     vl_logic_vector(7 downto 0);
        scb_bstsds_b    : in     vl_logic_vector(7 downto 0);
        scb_bstsds_c    : in     vl_logic_vector(7 downto 0);
        ffc_ck_core_tx  : in     vl_logic;
        ffc_ck_core_rx  : in     vl_logic;
        ffc_quad_rst    : in     vl_logic;
        ffc_macro_rst   : in     vl_logic;
        ffc_lane_tx_rst0: in     vl_logic;
        ffc_lane_tx_rst1: in     vl_logic;
        ffc_lane_tx_rst2: in     vl_logic;
        ffc_lane_tx_rst3: in     vl_logic;
        ffc_lane_rx_rst0: in     vl_logic;
        ffc_lane_rx_rst1: in     vl_logic;
        ffc_lane_rx_rst2: in     vl_logic;
        ffc_lane_rx_rst3: in     vl_logic;
        ffc_pcie_ei_en_0: in     vl_logic;
        ffc_pcie_ei_en_1: in     vl_logic;
        ffc_pcie_ei_en_2: in     vl_logic;
        ffc_pcie_ei_en_3: in     vl_logic;
        ffc_pcie_ct_0   : in     vl_logic;
        ffc_pcie_ct_1   : in     vl_logic;
        ffc_pcie_ct_2   : in     vl_logic;
        ffc_pcie_ct_3   : in     vl_logic;
        ffs_pcie_con_0  : out    vl_logic;
        ffs_pcie_con_1  : out    vl_logic;
        ffs_pcie_con_2  : out    vl_logic;
        ffs_pcie_con_3  : out    vl_logic;
        ffs_pcie_done_0 : out    vl_logic;
        ffs_pcie_done_1 : out    vl_logic;
        ffs_pcie_done_2 : out    vl_logic;
        ffs_pcie_done_3 : out    vl_logic;
        ffc_pcie_tx_0   : in     vl_logic;
        ffc_pcie_tx_1   : in     vl_logic;
        ffc_pcie_tx_2   : in     vl_logic;
        ffc_pcie_tx_3   : in     vl_logic;
        ffc_pcie_rx_0   : in     vl_logic;
        ffc_pcie_rx_1   : in     vl_logic;
        ffc_pcie_rx_2   : in     vl_logic;
        ffc_pcie_rx_3   : in     vl_logic;
        ffc_sd_0        : in     vl_logic;
        ffc_sd_1        : in     vl_logic;
        ffc_sd_2        : in     vl_logic;
        ffc_sd_3        : in     vl_logic;
        ffc_en_cga_0    : in     vl_logic;
        ffc_en_cga_1    : in     vl_logic;
        ffc_en_cga_2    : in     vl_logic;
        ffc_en_cga_3    : in     vl_logic;
        ffc_align_en_0  : in     vl_logic;
        ffc_align_en_1  : in     vl_logic;
        ffc_align_en_2  : in     vl_logic;
        ffc_align_en_3  : in     vl_logic;
        ffc_ab_reset    : in     vl_logic;
        ffc_cd_reset    : in     vl_logic;
        ffs_ls_status_0 : out    vl_logic;
        ffs_ls_status_1 : out    vl_logic;
        ffs_ls_status_2 : out    vl_logic;
        ffs_ls_status_3 : out    vl_logic;
        ffs_ab_status   : out    vl_logic;
        ffs_cd_status   : out    vl_logic;
        ffs_ab_aligned  : out    vl_logic;
        ffs_cd_aligned  : out    vl_logic;
        ffs_ab_failed   : out    vl_logic;
        ffs_cd_failed   : out    vl_logic;
        ffc_fb_lb_0     : in     vl_logic;
        ffc_fb_lb_1     : in     vl_logic;
        ffc_fb_lb_2     : in     vl_logic;
        ffc_fb_lb_3     : in     vl_logic;
        ffc_sb_inv_rx_0 : in     vl_logic;
        ffc_sb_inv_rx_1 : in     vl_logic;
        ffc_sb_inv_rx_2 : in     vl_logic;
        ffc_sb_inv_rx_3 : in     vl_logic;
        ffs_cc_orun_0   : out    vl_logic;
        ffs_cc_orun_1   : out    vl_logic;
        ffs_cc_orun_2   : out    vl_logic;
        ffs_cc_orun_3   : out    vl_logic;
        ffs_cc_urun_0   : out    vl_logic;
        ffs_cc_urun_1   : out    vl_logic;
        ffs_cc_urun_2   : out    vl_logic;
        ffs_cc_urun_3   : out    vl_logic;
        addro           : out    vl_logic_vector(7 downto 0);
        wdatao          : out    vl_logic_vector(7 downto 0);
        rdo             : out    vl_logic;
        wstbo           : out    vl_logic;
        rdatai          : in     vl_logic_vector(7 downto 0);
        inti            : in     vl_logic;
        rdatao          : out    vl_logic_vector(7 downto 0);
        into            : out    vl_logic;
        addri           : in     vl_logic_vector(7 downto 0);
        wdatai          : in     vl_logic_vector(7 downto 0);
        rdi             : in     vl_logic;
        wstbi           : in     vl_logic;
        cs_chif_0       : in     vl_logic;
        cs_chif_1       : in     vl_logic;
        cs_chif_2       : in     vl_logic;
        cs_chif_3       : in     vl_logic;
        cs_qif          : in     vl_logic;
        pwrupres        : in     vl_logic;
        testclk         : out    vl_logic;
        testclk_maco    : in     vl_logic;
        ff_sysclk_p1    : out    vl_logic;
        ff_sysclk0      : out    vl_logic;
        ff_sysclk1      : out    vl_logic;
        ff_sysclk2      : out    vl_logic;
        ff_sysclk3      : out    vl_logic;
        ff_rxclk_p1     : out    vl_logic;
        ff_rxclk_p2     : out    vl_logic;
        ff_rxclk0       : out    vl_logic;
        ff_rxclk1       : out    vl_logic;
        ff_rxclk2       : out    vl_logic;
        ff_rxclk3       : out    vl_logic;
        quad_clk        : out    vl_logic;
        grp_clk_p1      : in     vl_logic_vector(3 downto 0);
        grp_clk_p2      : in     vl_logic_vector(3 downto 0);
        grp_start       : in     vl_logic_vector(3 downto 0);
        grp_done        : in     vl_logic_vector(3 downto 0);
        grp_deskew_error: in     vl_logic_vector(3 downto 0);
        iqa_start_ls    : out    vl_logic;
        iqa_done_ls     : out    vl_logic;
        iqa_and_fp1_ls  : out    vl_logic;
        iqa_and_fp0_ls  : out    vl_logic;
        iqa_or_fp1_ls   : out    vl_logic;
        iqa_or_fp0_ls   : out    vl_logic;
        iqa_rst_n       : out    vl_logic;
        ff_tclk0        : in     vl_logic;
        ff_tclk1        : in     vl_logic;
        ff_tclk2        : in     vl_logic;
        ff_tclk3        : in     vl_logic;
        ff_rclk0        : in     vl_logic;
        ff_rclk1        : in     vl_logic;
        ff_rclk2        : in     vl_logic;
        ff_rclk3        : in     vl_logic;
        ff_txd_0        : in     vl_logic_vector(23 downto 0);
        fb_rxd_0        : out    vl_logic_vector(23 downto 0);
        ff_txd_1        : in     vl_logic_vector(23 downto 0);
        fb_rxd_1        : out    vl_logic_vector(23 downto 0);
        ff_txd_2        : in     vl_logic_vector(23 downto 0);
        fb_rxd_2        : out    vl_logic_vector(23 downto 0);
        ff_txd_3        : in     vl_logic_vector(23 downto 0);
        fb_rxd_3        : out    vl_logic_vector(23 downto 0);
        cout            : out    vl_logic_vector(21 downto 0);
        serdes_cout     : out    vl_logic_vector(21 downto 0);
        tck_fmac        : out    vl_logic;
        tck_fmacp       : in     vl_logic;
        cin             : in     vl_logic_vector(12 downto 0);
        serdes_coutp    : in     vl_logic_vector(21 downto 0);
        coutp           : in     vl_logic_vector(21 downto 0);
        quad_id         : in     vl_logic_vector(1 downto 0);
        bs2pad_0        : in     vl_logic;
        bs2pad_1        : in     vl_logic;
        bs2pad_2        : in     vl_logic;
        bs2pad_3        : in     vl_logic;
        bs_tx_sel       : in     vl_logic;
        bs_rx_ref_sel   : in     vl_logic;
        bs4pad_0        : out    vl_logic;
        bs4pad_1        : out    vl_logic;
        bs4pad_2        : out    vl_logic;
        bs4pad_3        : out    vl_logic;
        bs4refck        : out    vl_logic;
        bs4rxrefck      : out    vl_logic;
        grp0_wrst_in_n  : in     vl_logic;
        grp1_wrst_in_n  : in     vl_logic;
        grp2_wrst_in_n  : in     vl_logic;
        grp3_wrst_in_n  : in     vl_logic;
        grp0_rrst_in_n  : in     vl_logic;
        grp1_rrst_in_n  : in     vl_logic;
        grp2_rrst_in_n  : in     vl_logic;
        grp3_rrst_in_n  : in     vl_logic;
        is_slave0_in    : in     vl_logic;
        is_slave1_in    : in     vl_logic;
        is_slave2_in    : in     vl_logic;
        is_slave3_in    : in     vl_logic;
        grp0_wrst_Lout_n: out    vl_logic;
        grp1_wrst_Lout_n: out    vl_logic;
        grp2_wrst_Lout_n: out    vl_logic;
        grp3_wrst_Lout_n: out    vl_logic;
        grp0_rrst_Lout_n: out    vl_logic;
        grp1_rrst_Lout_n: out    vl_logic;
        grp2_rrst_Lout_n: out    vl_logic;
        grp3_rrst_Lout_n: out    vl_logic;
        is_slave0_Lout  : out    vl_logic;
        is_slave1_Lout  : out    vl_logic;
        is_slave2_Lout  : out    vl_logic;
        is_slave3_Lout  : out    vl_logic;
        grp0_wrst_Rout_n: out    vl_logic;
        grp1_wrst_Rout_n: out    vl_logic;
        grp2_wrst_Rout_n: out    vl_logic;
        grp3_wrst_Rout_n: out    vl_logic;
        grp0_rrst_Rout_n: out    vl_logic;
        grp1_rrst_Rout_n: out    vl_logic;
        grp2_rrst_Rout_n: out    vl_logic;
        grp3_rrst_Rout_n: out    vl_logic;
        is_slave0_Rout  : out    vl_logic;
        is_slave1_Rout  : out    vl_logic;
        is_slave2_Rout  : out    vl_logic;
        is_slave3_Rout  : out    vl_logic;
        TIE_HIGH        : out    vl_logic;
        TIE_LOW         : out    vl_logic;
        ffs_rlos_lo0    : out    vl_logic;
        ffs_rlos_lo1    : out    vl_logic;
        ffs_rlos_lo2    : out    vl_logic;
        ffs_rlos_lo3    : out    vl_logic
    );
end pcs_quad_top;
