library verilog;
use verilog.vl_types.all;
entity e2top_quad is
    port(
        ECP2M_35K       : in     vl_logic;
        HDINP0          : in     vl_logic;
        HDINN0          : in     vl_logic;
        HDINP1          : in     vl_logic;
        HDINN1          : in     vl_logic;
        HDINP2          : in     vl_logic;
        HDINN2          : in     vl_logic;
        HDINP3          : in     vl_logic;
        HDINN3          : in     vl_logic;
        sync_pulse      : in     vl_logic;
        REFCLKP         : in     vl_logic;
        REFCLKN         : in     vl_logic;
        ck_core_tx      : in     vl_logic;
        ck_core_rx      : in     vl_logic;
        macrorst        : in     vl_logic;
        macropdb        : in     vl_logic;
        pwr_on_rst      : in     vl_logic;
        rrst            : in     vl_logic_vector(3 downto 0);
        trst            : in     vl_logic;
        td0             : in     vl_logic_vector(9 downto 0);
        td1             : in     vl_logic_vector(9 downto 0);
        td2             : in     vl_logic_vector(9 downto 0);
        td3             : in     vl_logic_vector(9 downto 0);
        bs2pad_0        : in     vl_logic;
        bs2pad_1        : in     vl_logic;
        bs2pad_2        : in     vl_logic;
        bs2pad_3        : in     vl_logic;
        rx_bs_mode      : in     vl_logic;
        tx_bs_mode      : in     vl_logic;
        pcie_mode       : in     vl_logic;
        pci_det_ct0     : in     vl_logic;
        pci_det_ct1     : in     vl_logic;
        pci_det_ct2     : in     vl_logic;
        pci_det_ct3     : in     vl_logic;
        pci_det_en0     : in     vl_logic;
        pci_det_en1     : in     vl_logic;
        pci_det_en2     : in     vl_logic;
        pci_det_en3     : in     vl_logic;
        pci_ei_en0      : in     vl_logic;
        pci_ei_en1      : in     vl_logic;
        pci_ei_en2      : in     vl_logic;
        pci_ei_en3      : in     vl_logic;
        ser_ctl_qd_0    : in     vl_logic_vector(7 downto 0);
        ser_ctl_qd_1    : in     vl_logic_vector(7 downto 0);
        ser_ctl_qd_2    : in     vl_logic_vector(7 downto 0);
        ser_ctl_qd_3    : in     vl_logic_vector(7 downto 0);
        ser_ctl_qd_4    : in     vl_logic_vector(7 downto 0);
        ser_ctl_ch0_0   : in     vl_logic_vector(7 downto 0);
        ser_ctl_ch0_1   : in     vl_logic_vector(7 downto 0);
        ser_ctl_ch0_2   : in     vl_logic_vector(7 downto 0);
        ser_ctl_ch0_3   : in     vl_logic_vector(7 downto 0);
        ser_ctl_ch0_4   : in     vl_logic_vector(7 downto 0);
        ser_ctl_ch1_0   : in     vl_logic_vector(7 downto 0);
        ser_ctl_ch1_1   : in     vl_logic_vector(7 downto 0);
        ser_ctl_ch1_2   : in     vl_logic_vector(7 downto 0);
        ser_ctl_ch1_3   : in     vl_logic_vector(7 downto 0);
        ser_ctl_ch1_4   : in     vl_logic_vector(7 downto 0);
        ser_ctl_ch2_0   : in     vl_logic_vector(7 downto 0);
        ser_ctl_ch2_1   : in     vl_logic_vector(7 downto 0);
        ser_ctl_ch2_2   : in     vl_logic_vector(7 downto 0);
        ser_ctl_ch2_3   : in     vl_logic_vector(7 downto 0);
        ser_ctl_ch2_4   : in     vl_logic_vector(7 downto 0);
        ser_ctl_ch3_0   : in     vl_logic_vector(7 downto 0);
        ser_ctl_ch3_1   : in     vl_logic_vector(7 downto 0);
        ser_ctl_ch3_2   : in     vl_logic_vector(7 downto 0);
        ser_ctl_ch3_3   : in     vl_logic_vector(7 downto 0);
        ser_ctl_ch3_4   : in     vl_logic_vector(7 downto 0);
        ser_mem_ch0     : in     vl_logic_vector(81 downto 0);
        ser_mem_ch1     : in     vl_logic_vector(81 downto 0);
        ser_mem_ch2     : in     vl_logic_vector(81 downto 0);
        ser_mem_ch3     : in     vl_logic_vector(81 downto 0);
        ser_mem_qd      : in     vl_logic_vector(71 downto 0);
        VCCIB0          : in     vl_logic;
        VCCIB1          : in     vl_logic;
        VCCIB2          : in     vl_logic;
        VCCIB3          : in     vl_logic;
        VCCOB0          : in     vl_logic;
        VCCOB1          : in     vl_logic;
        VCCOB2          : in     vl_logic;
        VCCOB3          : in     vl_logic;
        VCCAX33         : in     vl_logic;
        VCCRX0          : in     vl_logic;
        VCCRX1          : in     vl_logic;
        VCCRX2          : in     vl_logic;
        VCCRX3          : in     vl_logic;
        VCCTX0          : in     vl_logic;
        VCCTX1          : in     vl_logic;
        VCCTX2          : in     vl_logic;
        VCCTX3          : in     vl_logic;
        VCCP            : in     vl_logic;
        VSSQ            : in     vl_logic;
        HDOUTP0         : out    vl_logic;
        HDOUTN0         : out    vl_logic;
        HDOUTP1         : out    vl_logic;
        HDOUTN1         : out    vl_logic;
        HDOUTP2         : out    vl_logic;
        HDOUTN2         : out    vl_logic;
        HDOUTP3         : out    vl_logic;
        HDOUTN3         : out    vl_logic;
        rd0             : out    vl_logic_vector(9 downto 0);
        rd1             : out    vl_logic_vector(9 downto 0);
        rd2             : out    vl_logic_vector(9 downto 0);
        rd3             : out    vl_logic_vector(9 downto 0);
        rck0            : out    vl_logic;
        rck1            : out    vl_logic;
        rck2            : out    vl_logic;
        rck3            : out    vl_logic;
        tck0            : out    vl_logic;
        tck1            : out    vl_logic;
        tck2            : out    vl_logic;
        tck3            : out    vl_logic;
        pci_connect0    : out    vl_logic;
        pci_connect1    : out    vl_logic;
        pci_connect2    : out    vl_logic;
        pci_connect3    : out    vl_logic;
        pci_det_done0   : out    vl_logic;
        pci_det_done1   : out    vl_logic;
        pci_det_done2   : out    vl_logic;
        pci_det_done3   : out    vl_logic;
        plol            : out    vl_logic;
        rlol            : out    vl_logic_vector(3 downto 0);
        rlos_hi         : out    vl_logic_vector(3 downto 0);
        rlos_lo         : out    vl_logic_vector(3 downto 0);
        ser_sts_qd_0    : out    vl_logic_vector(7 downto 0);
        ser_sts_qd_1    : out    vl_logic_vector(7 downto 0);
        ser_sts_ch0_1   : out    vl_logic_vector(7 downto 0);
        ser_sts_ch0_2   : out    vl_logic_vector(7 downto 0);
        ser_sts_ch0_3   : out    vl_logic_vector(7 downto 0);
        ser_sts_ch1_1   : out    vl_logic_vector(7 downto 0);
        ser_sts_ch1_2   : out    vl_logic_vector(7 downto 0);
        ser_sts_ch1_3   : out    vl_logic_vector(7 downto 0);
        ser_sts_ch2_1   : out    vl_logic_vector(7 downto 0);
        ser_sts_ch2_2   : out    vl_logic_vector(7 downto 0);
        ser_sts_ch2_3   : out    vl_logic_vector(7 downto 0);
        ser_sts_ch3_1   : out    vl_logic_vector(7 downto 0);
        ser_sts_ch3_2   : out    vl_logic_vector(7 downto 0);
        ser_sts_ch3_3   : out    vl_logic_vector(7 downto 0);
        refck2core      : out    vl_logic;
        tck_full        : out    vl_logic;
        oob_out0        : out    vl_logic;
        oob_out1        : out    vl_logic;
        oob_out2        : out    vl_logic;
        oob_out3        : out    vl_logic;
        bs4pad_0        : out    vl_logic;
        bs4pad_1        : out    vl_logic;
        bs4pad_2        : out    vl_logic;
        bs4pad_3        : out    vl_logic;
        bs4refck        : out    vl_logic
    );
end e2top_quad;
