-- $Header: //synplicity/map202003lat/mappers/cpld/lib/gen_mach/add.vhd#1 $
@ER--qC88sFRl8CkDRsVFRb#kCFsOFDD5NH00OHCR#qbvBj]6jXjv2H
DLssN$ RQ 
 ;kR#CQ   38#0_oDFH4O_43ncN;DD
M
C0$H0R7q7R
H#
MoCCOsH58IH0:ERR0HMCsoC:.=4U
2;
sbF0
5
qR,A:MRHR8#0_oDFHPO_CFO0sH5I8-0E4FR8IFM0R;j2
R
RRRRRRQRBhH:RM0R#8F_Do;HO
R
m:kRF00R#8F_Do_HOP0COFIs5HE80-84RF0IMF2Rj;B

mRza:kRF00R#8F_Do
HO

2;
8CMR7q7;N

sHOE00COkRsCpqe_7F7RV7Rq7#RH
F
OlMbFCRM0B_Bzq
77RbRRF5s0
RRRRqRRjRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR:RRHMR1RRap7_mBtQ;R
RRRRRARjRRRRRRRRRRRRRRRRRRRRRRRRRR:RRRMRHRRRR1_a7pQmtBR;
RRRRRhBQRRRRRRRRRRRRRRRRRRRRRRRRRRRR:HRRMRRRR71a_tpmQ
B;RRRRRjR1RRRRRRRRRRRRRRRRRRRRRRRRRRRRRR:RFRk0RaR17m_pt;QB
RRRRBRRmRzaRRRRRRRRRRRRRRRRRRRRRRRRRRR:R0FkR1RRap7_mBtQ2C;
MO8RFFlbM0CM;#

HNoMDNROsRs$RRR:#_08DHFoOC_POs0F5HRI8-0E4FR8IFM0R2jR;H
#oDMNRMOF#40_R#:R0D8_FOoH;L

CMoH
4Sz:BRBz7_q7mRu)vaRqRu5q25j,5RAjR2,B,QhRjm52O,RN$ss52j2;R
RRRRRR.Rp:FRVsRRHH4MRRR0FI0H8ER-4oCCMsCN0
RRRRRRRRRRRRRRRRRz.:BRBz7_q7mRu)vaRqRu5q25H,5RAHR2,OsNs$-5H4R2,m25H,NROs5s$H;22
RRRRRRRR8CMRMoCC0sNCR;
RRRRRBRRmRza<O=RN$ss5HRI8-0E4;R2
C

Mp8Re7_q7
;

