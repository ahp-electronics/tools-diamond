library verilog;
use verilog.vl_types.all;
entity njtag_qual is
    port(
        isc_data_shift_cq: out    vl_logic;
        isc_addr_shift_cq: out    vl_logic;
        verify_id_cq    : out    vl_logic;
        idcode_pub_cq   : out    vl_logic;
        uidcode_pub_cq  : out    vl_logic;
        usercode_cq     : out    vl_logic;
        usercode_dryrun_cq: out    vl_logic;
        prog_dryrun_addr_cq: out    vl_logic;
        read_temp_cq    : out    vl_logic;
        lsc_device_ctrl_cq: out    vl_logic;
        lsc_shift_password_cq: out    vl_logic;
        lsc_read_status_cq: out    vl_logic;
        lsc_read_status1_cq: out    vl_logic;
        lsc_check_busy_cq: out    vl_logic;
        lsc_refresh_cq  : out    vl_logic;
        lsc_bitstream_burst_cq: out    vl_logic;
        idcode_prv_cq   : out    vl_logic;
        lsc_read_pes_cq : out    vl_logic;
        lsc_prog_ctrl0_cq: out    vl_logic;
        lsc_read_ctrl0_cq: out    vl_logic;
        lsc_prog_ctrl1_cq: out    vl_logic;
        lsc_read_ctrl1_cq: out    vl_logic;
        lsc_reset_crc_cq: out    vl_logic;
        lsc_read_crc_cq : out    vl_logic;
        lsc_write_comp_dic_cq: out    vl_logic;
        sf_prog_ucode_cq: out    vl_logic;
        sf_program_cq   : out    vl_logic;
        sf_read_cq      : out    vl_logic;
        sf_erase_cq     : out    vl_logic;
        sf_prog_done_cq : out    vl_logic;
        sf_erase_done_cq: out    vl_logic;
        sf_prog_sec_cq  : out    vl_logic;
        sf_init_addr_cq : out    vl_logic;
        sf_write_addr_cq: out    vl_logic;
        sf_prog_incr_rti_cq: out    vl_logic;
        sf_prog_incr_enc_cq: out    vl_logic;
        sf_prog_incr_cmp_cq: out    vl_logic;
        sf_prog_incr_cne_cq: out    vl_logic;
        sf_vfy_incr_rti_cq: out    vl_logic;
        sf_prog_sed_crc_cq: out    vl_logic;
        sf_read_sed_crc_cq: out    vl_logic;
        sf_write_bus_addr_cq: out    vl_logic;
        sf_pcs_write_cq : out    vl_logic;
        sf_pcs_read_cq  : out    vl_logic;
        sf_ebr_write_cq : out    vl_logic;
        sf_ebr_read_cq  : out    vl_logic;
        fl_prog_ucode_cq: out    vl_logic;
        fl_erase_cq     : out    vl_logic;
        fl_prog_done_cq : out    vl_logic;
        fl_prog_sec_cq  : out    vl_logic;
        fl_prog_secplus_cq: out    vl_logic;
        fl_init_addr_cq : out    vl_logic;
        fl_write_addr_cq: out    vl_logic;
        fl_prog_incr_nv_cq: out    vl_logic;
        fl_read_incr_nv_cq: out    vl_logic;
        fl_prog_password_cq: out    vl_logic;
        fl_read_password_cq: out    vl_logic;
        fl_prog_cipher_key0_cq: out    vl_logic;
        fl_prog_cipher_key1_cq: out    vl_logic;
        fl_read_cipher_key0_cq: out    vl_logic;
        fl_read_cipher_key1_cq: out    vl_logic;
        fl_prog_feature_cq: out    vl_logic;
        fl_read_feature_cq: out    vl_logic;
        fl_prog_feabits_cq: out    vl_logic;
        fl_read_feabits_cq: out    vl_logic;
        fl_init_addr_ufm_cq: out    vl_logic;
        fl_prog_tag_cq  : out    vl_logic;
        fl_erase_tag_cq : out    vl_logic;
        fl_read_tag_cq  : out    vl_logic;
        fl_prog_csec_cq : out    vl_logic;
        fl_read_csec_cq : out    vl_logic;
        fl_prog_usec_cq : out    vl_logic;
        fl_read_usec_cq : out    vl_logic;
        fl_prog_authdone_cq: out    vl_logic;
        fl_prog_authmode_cq: out    vl_logic;
        fl_prog_aesfea_cq: out    vl_logic;
        fl_read_authmode_cq: out    vl_logic;
        fl_read_aesfea_cq: out    vl_logic;
        lsc_jump_cq     : out    vl_logic;
        lsc_chip_select_cq: out    vl_logic;
        lsc_flow_through_cq: out    vl_logic;
        bypass_cq       : out    vl_logic;
        sed_init_addr_cq: out    vl_logic;
        sed_write_addr_cq: out    vl_logic;
        sed_prog_incr_rti_cq: out    vl_logic;
        sed_prog_incr_cmp_cq: out    vl_logic;
        sed_prog_sed_crc_cq: out    vl_logic;
        sed_prog_ctrl0_cq: out    vl_logic;
        sed_prog_ctrl1_cq: out    vl_logic;
        sed_write_comp_dic_cq: out    vl_logic;
        lsc_i2ci_crbr_wt_cq: out    vl_logic;
        lsc_i2ci_txdr_wt_cq: out    vl_logic;
        lsc_i2ci_rxdr_rd_cq: out    vl_logic;
        lsc_i2ci_sr_rd_cq: out    vl_logic;
        lsc_auth_ctrl_cq: out    vl_logic;
        fl_prog_pubkey0_cq: out    vl_logic;
        fl_prog_pubkey1_cq: out    vl_logic;
        fl_prog_pubkey2_cq: out    vl_logic;
        fl_prog_pubkey3_cq: out    vl_logic;
        fl_read_pubkey0_cq: out    vl_logic;
        fl_read_pubkey1_cq: out    vl_logic;
        fl_read_pubkey2_cq: out    vl_logic;
        fl_read_pubkey3_cq: out    vl_logic;
        lsc_verify_uid_cq: out    vl_logic;
        lsc_erase_all_cq: out    vl_logic;
        lsc_alter_sec_cq: out    vl_logic;
        lsc_alter_sram_sec_cq: out    vl_logic;
        lsc_alter_port_sec_cq: out    vl_logic;
        lsc_prog_uds_cq : out    vl_logic;
        isc_nj_enabled  : in     vl_logic;
        isc_nj_disable_completing: in     vl_logic;
        njaccess_sram   : in     vl_logic;
        njaccess_flash  : in     vl_logic;
        njaccess_tag    : in     vl_logic;
        njenable_tran   : in     vl_logic;
        ctrl_tran_edit  : in     vl_logic;
        jtag_active_smsync: in     vl_logic;
        jburst_inp      : in     vl_logic;
        dryrun_inp      : in     vl_logic;
        sed_active      : in     vl_logic;
        bypass_c        : in     vl_logic;
        verify_id_c     : in     vl_logic;
        idcode_pub_c    : in     vl_logic;
        uidcode_pub_c   : in     vl_logic;
        usercode_c      : in     vl_logic;
        usercode_dryrun_c: in     vl_logic;
        prog_dryrun_addr_c: in     vl_logic;
        read_temp_c     : in     vl_logic;
        lsc_device_ctrl_c: in     vl_logic;
        lsc_shift_password_c: in     vl_logic;
        lsc_read_status_c: in     vl_logic;
        lsc_read_status1_c: in     vl_logic;
        lsc_check_busy_c: in     vl_logic;
        lsc_refresh_c   : in     vl_logic;
        lsc_bitstream_burst_c: in     vl_logic;
        lsc_i2ci_crbr_wt_c: in     vl_logic;
        lsc_i2ci_txdr_wt_c: in     vl_logic;
        lsc_i2ci_rxdr_rd_c: in     vl_logic;
        lsc_i2ci_sr_rd_c: in     vl_logic;
        idcode_prv_c    : in     vl_logic;
        read_pes_c      : in     vl_logic;
        isc_program_c   : in     vl_logic;
        isc_prog_ucode_c: in     vl_logic;
        isc_read_c      : in     vl_logic;
        isc_erase_c     : in     vl_logic;
        isc_prog_done_c : in     vl_logic;
        isc_erase_done_c: in     vl_logic;
        isc_prog_sec_c  : in     vl_logic;
        isc_prog_secplus_c: in     vl_logic;
        isc_data_shift_c: in     vl_logic;
        isc_addr_shift_c: in     vl_logic;
        lsc_init_addr_c : in     vl_logic;
        lsc_write_addr_c: in     vl_logic;
        lsc_prog_incr_rti_c: in     vl_logic;
        lsc_prog_incr_enc_c: in     vl_logic;
        lsc_prog_incr_cmp_c: in     vl_logic;
        lsc_prog_incr_cne_c: in     vl_logic;
        lsc_vfy_incr_rti_c: in     vl_logic;
        lsc_prog_ctrl0_c: in     vl_logic;
        lsc_read_ctrl0_c: in     vl_logic;
        lsc_prog_ctrl1_c: in     vl_logic;
        lsc_read_ctrl1_c: in     vl_logic;
        lsc_reset_crc_c : in     vl_logic;
        lsc_read_crc_c  : in     vl_logic;
        lsc_prog_sed_crc_c: in     vl_logic;
        lsc_read_sed_crc_c: in     vl_logic;
        lsc_prog_password_c: in     vl_logic;
        lsc_read_password_c: in     vl_logic;
        lsc_prog_cipher_key0_c: in     vl_logic;
        lsc_prog_cipher_key1_c: in     vl_logic;
        lsc_read_cipher_key0_c: in     vl_logic;
        lsc_read_cipher_key1_c: in     vl_logic;
        lsc_prog_feature_c: in     vl_logic;
        lsc_read_feature_c: in     vl_logic;
        lsc_prog_feabits_c: in     vl_logic;
        lsc_read_feabits_c: in     vl_logic;
        lsc_write_comp_dic_c: in     vl_logic;
        lsc_write_bus_addr_c: in     vl_logic;
        lsc_pcs_write_c : in     vl_logic;
        lsc_pcs_read_c  : in     vl_logic;
        lsc_ebr_write_c : in     vl_logic;
        lsc_ebr_read_c  : in     vl_logic;
        lsc_prog_incr_nv_c: in     vl_logic;
        lsc_read_incr_nv_c: in     vl_logic;
        lsc_init_addr_ufm_c: in     vl_logic;
        lsc_prog_tag_c  : in     vl_logic;
        lsc_erase_tag_c : in     vl_logic;
        lsc_read_tag_c  : in     vl_logic;
        lsc_prog_csec_c : in     vl_logic;
        lsc_read_csec_c : in     vl_logic;
        lsc_prog_usec_c : in     vl_logic;
        lsc_read_usec_c : in     vl_logic;
        lsc_prog_authdone_c: in     vl_logic;
        lsc_prog_authmode_c: in     vl_logic;
        lsc_prog_aesfea_c: in     vl_logic;
        lsc_read_authmode_c: in     vl_logic;
        lsc_read_aesfea_c: in     vl_logic;
        lsc_chip_select_c: in     vl_logic;
        lsc_flow_through_c: in     vl_logic;
        lsc_jump_c      : in     vl_logic;
        lsc_verify_uid_c: in     vl_logic;
        lsc_erase_all_c : in     vl_logic;
        lsc_auth_ctrl_c : in     vl_logic;
        lsc_prog_ecdsa_pubkey0_c: in     vl_logic;
        lsc_prog_ecdsa_pubkey1_c: in     vl_logic;
        lsc_prog_ecdsa_pubkey2_c: in     vl_logic;
        lsc_prog_ecdsa_pubkey3_c: in     vl_logic;
        lsc_read_ecdsa_pubkey0_c: in     vl_logic;
        lsc_read_ecdsa_pubkey1_c: in     vl_logic;
        lsc_read_ecdsa_pubkey2_c: in     vl_logic;
        lsc_read_ecdsa_pubkey3_c: in     vl_logic;
        lsc_alter_sec_c : in     vl_logic;
        lsc_alter_sram_sec_c: in     vl_logic;
        lsc_alter_port_sec_c: in     vl_logic;
        lsc_prog_uds_c  : in     vl_logic
    );
end njtag_qual;
