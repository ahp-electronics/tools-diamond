--
@ER--RbBF$osHE50RO42RgRgg1b$MDHHO0R$,Q3MO
R--RDqDRosHER0#sCC#s8PC3-
-

---f-R]8CNCRs:/$/#MHbDO$H0/blN.jj.jNdD0N/lbsbC#b/ODD8/HoL/CDM_NH00OOC/lDb_0E3P8Ry4f-
-
H
DLssN$CRHC
C;kR#CHCCC38#0_oDFH4O_43ncN;DD
Ck#RCHCC03#8F_Do_HON0sHED3NDC;
M00H$FROlsbNCO_NO_klLRH0HS#
b0Fs5S
SbRCJ:MRHR8#0_oDFH
O;SDSb0RR:H#MR0D8_FOoH;S
SDR0H:MRHR8#0_oDFH
O;SJSCHRR:H#MR0D8_FOoH;S
SD:0RR0FkR8#0_oDFH
O;SJSCRF:Rk#0R0D8_FOoH
;S2
8CMRlOFbCNs_ONOkLl_H
0;
ONsECH0Os0kCFRLFNDCMVRFRlOFbCNs_ONOkLl_HH0R#C
Lo
HMSRCJ<b=RCNJRMC8RJ
H;SRD0<b=RDI0RERCMCRJH=4R''DRC#DCR0
H;CRM8LDFFC;NM
-
-RONOkDlkNR0C0RECDs0RCD#k0sRVF0lREbCRsHCPFRk#DCCPDFROlsbNCD#
HNLssH$RC;CC
Ck#RCHCC03#8F_Do_HO4c4n3DND;#
kCCRHC#C30D8_FOoH_HNs0NE3D
D;CHM00O$RFNlbsNC_OlOkR
H#SMoCCOsHRS5
Sx#HCRR:HCM0o
CsS
2;SsbF0S5
SHD0RH:RM0R#8F_Do_HOP0COF#s5H-xC4FR8IFM0R;j2
CSSJ:HRRRHM#_08DHFoOC_POs0F5x#HCR-48MFI0jFR2S;
SRD0:kRF00R#8F_Do;HO
CSSJRR:FRk0#_08DHFoO2
S;M
C8FROlsbNCO_NO;kl
s
NO0EHCkO0sLCRFCFDNFMRVFROlsbNCO_NORklHS#
#MHoNDDRD:0RR8#0_oDFHPO_CFO0sH5#x8CRF0IMF2Rj;#
SHNoMDCRDJRR:#_08DHFoOC_POs0F5x#HCFR8IFM0R;j2
FSOlMbFCRM0ObFlN_sCNkOOlH_L0#RH
bSSF5s0
SSSbRCJ:MRHR8#0_oDFH
O;SbSSD:0RRRHM#_08DHFoOS;
S0SDHRR:H#MR0D8_FOoH;S
SSHCJRH:RM0R#8F_Do;HO
SSSD:0RR0FkR8#0_oDFH
O;SCSSJRR:FRk0#_08DHFoOS
S2S;
CRM8ObFlFMMC0L;
CMoHRD
SDj052=R<R''j;D
SCjJ52=R<R''4;p
S:FRVsRRMHjMRRR0F#CHx-o4RCsMCN
0CS:SORlOFbCNs_ONOkLl_Hb0RFRs0lRNb5S
SSJbCRR=>D5CJM
2,SCSSJ=HR>JRCH25M,S
SS0bDRR=>D5D0M
2,SDSS0=HR>0RDH25M,S
SSRCJ=D>RCMJ5+,42
SSSD=0R>DRD0+5M4S2
S
2;S8CMRMoCC0sNCS;
D<0R=DRD0H5#x;C2
JSCRR<=D5CJ#CHx2C;
ML8RFCFDN
M;
LDHs$NsRCHCCk;
#HCRC3CC#_08DHFoO4_4nNc3D
D;kR#CHCCC38#0_oDFHNO_sEH03DND;M
C0$H0RlOFbCNs_0LHR
H#SsbF0S5
S:NRRRHM#_08DHFoOS;
S:LRRRHM#_08DHFoOS;
SHD0RH:RM0R#8F_Do;HO
CSSJ:HRRRHM#_08DHFoOS;
SRD0:kRF00R#8F_Do;HO
CSSJRR:FRk0#_08DHFoO2
S;M
C8FROlsbNCH_L0
;
NEsOHO0C0CksRFLFDMCNRRFVObFlN_sCLRH0HL#
CMoHRC
SJ=R<RHCJR8NMR0MFRR5NGRFsL
2;SRD0<L=RRCIEMNR5RsGFRRL2=4R''DRC#DCR0
H;CRM8LDFFC;NM
H
DLssN$CRHC
C;kR#CHCCC38#0_oDFH4O_43ncN;DD
Ck#RCHCC03#8F_Do_HON0sHED3NDC;
M00H$FROlsbNC#RH
CSoMHCsO#R5HRxC:MRH0CCos;R2
FSbs50R
NSSRH:RM0R#8F_Do_HOP0COF#s5H-xC4FR8IFM0R;j2
LSSRH:RM0R#8F_Do_HOP0COF#s5H-xC4FR8IFM0R;j2
DSS0RR:FRk0#_08DHFoOS;
SRCJ:kRF00R#8F_Do
HOS
2;CRM8ObFlN;sC
s
NO0EHCkO0sLCRFCFDNFMRVFROlsbNC#RH
HS#oDMNR0bD,CRbJRR:#_08DHFoOC_POs0F5x#HCFR8IFM0R;j2
FSOlMbFCRM0ObFlN_sCLRH0HS#
SsbF0S5
SRSN:MRHR8#0_oDFH
O;SLSSRH:RM0R#8F_Do;HO
SSSDR0H:MRHR8#0_oDFH
O;SCSSJ:HRRRHM#_08DHFoOS;
S0SDRF:Rk#0R0D8_FOoH;S
SSRCJ:kRF00R#8F_Do
HOS;S2
MSC8FROlMbFC;M0
oLCHSM
b5CJj<2R=4R''S;
b5D0j<2R=jR''S;
tV:RFMsRRRHMjFR0Rx#HCR-4oCCMsCN0RS
SOO:RFNlbsLC_H
0RSbSSFRs0lRNb5S
SS=SN>MN52
,RSSSSLL=>5,M2RS
SS0SDHb=>DM052
,RSSSSC=JH>JbC5,M2RS
SS0SD=D>b0+5M4R2,
SSSS=CJ>JbC54M+2S
SS
2;S8CMRMoCC0sNCS;
D<0R=DRb0H5#x;C2
JSCRR<=b5CJ#CHx2C;
ML8RFCFDN
M;
LDHs$NsRCHCCk;
#HCRC3CC#_08DHFoO4_4nNc3D
D;kR#CHCCC38#0_oDFHNO_sEH03DND;M
C0$H0RuBv_RpaHR#
RoRRCsMCHIO5HE80RH:RMo0CC:sR=jRU2-;R-NR[oR
RRFRbsq05:MRHR8#0_oDFHPO_CFO0sH5I8R0E-84RF0IMF2Rj;R
RRRRRRARR:MRHR8#0_oDFHPO_CFO0sH5I8R0E-84RF0IMF2Rj;R
RRRRRRpRRaRR:FRk0#_08DHFoO
2;CRM8B_vup
a;
ONsECH0Os0kCFRLFNDCMVRFRbOl_RD0HS#
VOkM0MHFRDONO0OMRF5OMN#0M#0RxD,RC#NVxRR:HCM0o2CsR0sCkRsMHCM0oRCsHS#
PHNsNCLDRNDCVb0l,MsO0RR:HCM0o;Cs
CSLo
HMSCSDNlV0b=R:RR#x/CRDNxV#;S
SH5VR5R#xlRF8DVCN#Rx2=2RjRC0EMS
SSMsO0=R:RNDCVb0lRS;
S#CDCSR
SOSsM:0R=DR5C0NVl+bRR;42
CSSMH8RVS;
S0sCkRsMs0OM;C
SMO8RNODOM
0;
FSOMN#0Mv0RqvXBuRR:HCM0oRCs:c=R;O
SF0M#NRM0DVCN#CHxRH:RMo0CC:sR=qRvXuBv;O
SF0M#NRM0OOlbM:0RR0HMCsoCRR:=OONDO5M0I0H8EC,DNHV#x;C2
SS
VOkM0MHFRGlNLRH05MOF#M0N0RRM:MRH0CCoss2RCs0kMMRH0CCos#RH
NSPsLHNDlCRN:GRR0HMCsoC;L
SCMoH
lSSN:GR=MR5+*42DVCN#CHxR4-R;S
SH5VRlRNG>I=RHE802ER0CSM
SNSlG=R:R8IH04E-;S
SCRM8H
V;SCSs0MksRGlN;C
SMl8RNHGL0
;
So#HMRNDoRD0:0R#8F_Do_HOP0COFOs5lMbO0R-48MFI0jFR2S;
#MHoNoDRC:JRR8#0_oDFHPO_CFO0sl5Ob0OM-84RF0IMF2Rj;S

ObFlFMMC0FROlsbNC#RH
oSSCsMCH5OR#CHxRH:RMo0CC;s2
bSSFRs05S
SS:NRRRHM#_08DHFoOC_POs0F5x#HCR-48MFI0jFR2S;
SRSL:MRHR8#0_oDFHPO_CFO0sH5#x4C-RI8FMR0Fj
2;SDSS0RR:FRk0#_08DHFoOS;
SJSCRF:Rk#0R0D8_FOoH
2SS;C
SMO8RFFlbM0CM;O
SFFlbM0CMRlOFbCNs_ONOkHlR#S
SoCCMsRHO5S
SSx#HCRR:HCM0o
CsS;S2
bSSF5s0
SSSDR0H:MRHR8#0_oDFHPO_CFO0sH5#x4C-RI8FMR0Fj
2;SCSSJ:HRRRHM#_08DHFoOC_POs0F5x#HCR-48MFI0jFR2S;
S0SDRF:Rk#0R0D8_FOoH;S
SSRCJ:kRF00R#8F_Do
HOS;S2
MSC8FROlMbFC;M0
#
SHNoMDJRCR#:R0D8_FOoH;L

CMoH
-S-RCk#R0NRIDF-CDPCRFDF	CNEN#8ROlECCA
S:VRHRH5I8R0E>qRvXuBv2CRoMNCs0
CRS:StRsVFRHMRMlROb0OM-84RF0IMFRRjoCCMsCN0
SSSO#FM00NMRLlG0RR:HCM0oRCs:l=RNHGL025M;S
SSMOF#M0N0MRlL:0RR0HMCsoCRR:=MC*DNHV#x
C;SCSLo
HMSBSS:FROlsbNCCRoMHCsONRlb#R5HRxC=4>R+LlG0M-lL
02SSSSb0FsRblNRS5
SSSSN>R=RlN5GRL08MFI0lFRM2L0,S
SSLSSRR=>LG5lL80RF0IMFMRlL,02
SSSS0SD=o>RDM052S,
SSSSC>J=RJoC5
M2SSSS2S;
S8CMRMoCC0sNC
;
S:SNRlOFbCNs_ONOk
lRSoSSCsMCHlORN5bR
SSSSx#HC>R=RbOlO
M0S2SS
SSSb0FsRblNRS5
SDSS0=HR>DRo0S,
SCSSJ=HR>CRoJS,
SDSS0>R=R,D0
SSSSRCJ=C>RJS
SS
2;S8CMRMoCC0sNC
;
SR--kR#CNHRsbCbDRlOFbCNs
:S1RRHV58IH0<ER=qRvXuBv2CRoMNCs0SC
SRB:ObFlNRsCoCCMsRHOlRNb5x#HCI=>HE802S
SSsbF0NRlb
R5SSSSN>R=R
N,SSSSL>R=R
L,SSSSD>0=R,D0
SSSS=CJ>JRC
SSS2S;
CRM8oCCMsCN0;C

ML8RFCFDN
M;
