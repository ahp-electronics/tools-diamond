--***************************************************************
-- 4-bit decade up counters with asynchronous clear, enable, and parallel data load.
-- -XiaoQiu ZHOU
--***************************************************************
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.std_logic_unsigned.ALL;
USE ieee.std_logic_arith.ALL;

ENTITY CDU14 IS 
    PORT (
        D0 : IN std_logic;
        D1 : IN std_logic;
        D2 : IN std_logic;
        D3 : IN std_logic;
        CLK : IN std_logic;
        LD : IN std_logic;
        EN : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic
    );
END CDU14;

ARCHITECTURE lattice_behav OF CDU14 IS
    SIGNAL Q_i  : std_logic_vector(3 downto 0);
BEGIN

PROCESS (CLK, LD, D0, D1, D2, D3, EN, CD)
BEGIN
  IF (CD = '1') THEN
    Q_i <= "0000";
  ELSIF rising_edge(CLK) THEN
    IF (LD = '1') THEN
      Q_i <= D3&D2&D1&D0;	
    ELSIF (EN = '1' AND (Q_i(3)='0' OR ( Q_i(2)='0' AND Q_i(1)='0' ))) THEN
      IF (Q_i = "1001") THEN
        Q_i <= "0000";	
      ELSE
        Q_i <= Q_i + 1;
	    END IF;  
	  END IF;  
  END IF;
end process;

Q0 <= Q_i(0);
Q1 <= Q_i(1);
Q2 <= Q_i(2);
Q3 <= Q_i(3);

END lattice_behav;
