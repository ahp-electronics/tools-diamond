library verilog;
use verilog.vl_types.all;
entity pcs_ch_dp is
    generic(
        TIE_LO_STS      : integer := 0
    );
    port(
        tx_clk          : in     vl_logic;
        rst_tx_clk_n    : in     vl_logic;
        rx_clk          : in     vl_logic;
        rst_rx_clk_n    : in     vl_logic;
        ebrd_clk        : in     vl_logic;
        rst_ebrd_clk_n  : in     vl_logic;
        fb_clk          : in     vl_logic;
        rst_fb_clk_n    : in     vl_logic;
        fft_clk         : in     vl_logic;
        ffr_clk         : in     vl_logic;
        txd_fifo_lb     : in     vl_logic_vector(9 downto 0);
        serdes_rxd      : in     vl_logic_vector(9 downto 0);
        sb_txd          : out    vl_logic_vector(9 downto 0);
        tobist_data     : out    vl_logic_vector(9 downto 0);
        bist_rx_data_sel: in     vl_logic;
        fmbist_data     : in     vl_logic_vector(9 downto 0);
        ff_tx_d         : in     vl_logic_vector(23 downto 0);
        ff_rx_d         : out    vl_logic_vector(23 downto 0);
        ffc_signal_detect: in     vl_logic;
        ffc_enable_cgalign: in     vl_logic;
        ffc_fb_loopback : in     vl_logic;
        ffc_sb_pfifo_lp : in     vl_logic;
        ffc_sb_inv_rx   : in     vl_logic;
        ffs_ls_sync_status: out    vl_logic;
        ffs_cc_overrun  : out    vl_logic;
        ffs_cc_underrun : out    vl_logic;
        ffs_rxfbfifo_error: out    vl_logic;
        ffs_txfbfifo_error: out    vl_logic;
        pcie_det_done   : in     vl_logic;
        pcie_connect    : in     vl_logic;
        pfifo_clr       : out    vl_logic;
        pfifo_clr_sel   : out    vl_logic;
        asyn_mode       : out    vl_logic;
        ffc_ei_en       : in     vl_logic;
        tsd_pcie_ei_en  : out    vl_logic;
        pcie_det_time_sel: out    vl_logic_vector(1 downto 0);
        sel_test_clk    : out    vl_logic;
        rx_ch           : out    vl_logic;
        bistrun_a1      : in     vl_logic;
        bistfc_a1       : in     vl_logic;
        bistdone_a1     : out    vl_logic_vector(1 downto 0);
        bistf_a1        : out    vl_logic_vector(1 downto 0);
        char_test_data  : in     vl_logic_vector(9 downto 0);
        char_test_mode  : in     vl_logic;
        pfifo_error     : in     vl_logic;
        prbs_error      : out    vl_logic;
        pcs_ctl_1_ch_00 : in     vl_logic_vector(7 downto 0);
        pcs_ctl_2_ch_01 : in     vl_logic_vector(7 downto 0);
        pcs_ctl_3_ch_02 : in     vl_logic_vector(7 downto 0);
        pcs_ctl_4_ch_03 : in     vl_logic_vector(7 downto 0);
        pcs_ctl_6_ch_05 : in     vl_logic_vector(7 downto 0);
        pcs_ctl_7_ch_06 : in     vl_logic_vector(7 downto 0);
        pcs_sts_1_ch_20 : out    vl_logic_vector(7 downto 0);
        pcs_sts_3_ch_22 : out    vl_logic_vector(7 downto 0);
        pcs_sts_5_ch_24 : out    vl_logic_vector(7 downto 0);
        pcs_sts_6_ch_25 : out    vl_logic_vector(7 downto 0);
        uc_mode         : in     vl_logic;
        fc_mode         : in     vl_logic;
        pcie_mode       : in     vl_logic;
        rio_mode        : in     vl_logic;
        xge_mode        : in     vl_logic;
        pcs_ctl_3_qd_02 : in     vl_logic_vector(7 downto 0);
        pcs_ctl_4_qd_03 : in     vl_logic_vector(7 downto 0);
        pcs_ctl_5_qd_04 : in     vl_logic_vector(7 downto 0);
        pcs_ctl_6_qd_05 : in     vl_logic_vector(7 downto 0);
        pcs_ctl_7_qd_06 : in     vl_logic_vector(7 downto 0);
        pcs_ctl_8_qd_07 : in     vl_logic_vector(7 downto 0);
        pcs_ctl_9_qd_08 : in     vl_logic_vector(7 downto 0);
        pcs_ctl_10_qd_09: in     vl_logic_vector(7 downto 0);
        pcs_ctl_11_qd_0a: in     vl_logic_vector(7 downto 0);
        pcs_ctl_12_qd_0b: in     vl_logic_vector(7 downto 0);
        pcs_ctl_13_qd_0c: in     vl_logic_vector(7 downto 0)
    );
end pcs_ch_dp;
