/* Because of the copyright that the IEEE has placed on IEEE 1801-2009 standard,
   Mentor Graphics cannot redistribute all the source code of this package to
   our customers.


   The missing source may be found in Annex B.2 of the IEEE 1801-2009 standard.*/
