library verilog;
use verilog.vl_types.all;
entity del1 is
    port(
        A               : in     vl_logic;
        Z               : out    vl_logic
    );
end del1;
