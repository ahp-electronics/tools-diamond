package mgc_rnm_pkg;
    nettype real wreal1driver with MGC_res_wreal1driver;
    nettype real wreal4state with MGC_res_wreal4state;
    nettype real wrealmin with MGC_res_wrealmin;
    nettype real wrealmax with MGC_res_wrealmax;
    nettype real wrealsum with MGC_res_wrealsum;
    nettype real wrealavg with MGC_res_wrealavg; 
endpackage

