library verilog;
use verilog.vl_types.all;
entity RS_UDP is
    -- This module cannot be connected to from
    -- VHDL because it has unnamed ports.
end RS_UDP;
