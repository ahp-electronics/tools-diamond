library verilog;
use verilog.vl_types.all;
entity pcs_quad is
    port(
        cin             : in     vl_logic_vector(11 downto 0);
        cyawstn         : in     vl_logic;
        ebrd_i_clk      : in     vl_logic_vector(3 downto 0);
        fb_i_clk        : in     vl_logic_vector(3 downto 0);
        ff_ebrd_clk     : in     vl_logic_vector(3 downto 0);
        ff_rxi_clk      : in     vl_logic_vector(3 downto 0);
        ff_tx_d_0       : in     vl_logic_vector(23 downto 0);
        ff_tx_d_1       : in     vl_logic_vector(23 downto 0);
        ff_tx_d_2       : in     vl_logic_vector(23 downto 0);
        ff_tx_d_3       : in     vl_logic_vector(23 downto 0);
        ff_txi_clk      : in     vl_logic_vector(3 downto 0);
        ffc_ei_en       : in     vl_logic_vector(3 downto 0);
        ffc_enable_cgalign: in     vl_logic_vector(3 downto 0);
        ffc_fb_loopback : in     vl_logic_vector(3 downto 0);
        ffc_lane_rx_rst : in     vl_logic_vector(3 downto 0);
        ffc_lane_tx_rst : in     vl_logic_vector(3 downto 0);
        ffc_macro_rst   : in     vl_logic;
        ffc_pci_det_en  : in     vl_logic_vector(3 downto 0);
        ffc_pcie_ct     : in     vl_logic_vector(3 downto 0);
        ffc_pfifo_clr   : in     vl_logic_vector(3 downto 0);
        ffc_quad_rst    : in     vl_logic;
        ffc_rrst        : in     vl_logic_vector(3 downto 0);
        ffc_rxpwdnb     : in     vl_logic_vector(3 downto 0);
        ffc_sb_inv_rx   : in     vl_logic_vector(3 downto 0);
        ffc_sb_pfifo_lp : in     vl_logic_vector(3 downto 0);
        ffc_signal_detect: in     vl_logic_vector(3 downto 0);
        ffc_sync_toggle : in     vl_logic;
        ffc_trst        : in     vl_logic;
        ffc_txpwdnb     : in     vl_logic_vector(3 downto 0);
        ffc_rx_div11_clk: in     vl_logic_vector(3 downto 0);
        ffc_tx_div11_clk: in     vl_logic_vector(3 downto 0);
        ffc_rx_rate_mode: in     vl_logic_vector(3 downto 0);
        ffc_tx_rate_mode: in     vl_logic_vector(3 downto 0);
        ffr_i_clk       : in     vl_logic_vector(3 downto 0);
        fft_i_clk       : in     vl_logic_vector(3 downto 0);
        ffc_ldr_core2tx_en: in     vl_logic_vector(3 downto 0);
        mc1_chif_ctl_ch0: in     vl_logic_vector(207 downto 0);
        mc1_chif_ctl_ch1: in     vl_logic_vector(207 downto 0);
        mc1_chif_ctl_ch2: in     vl_logic_vector(207 downto 0);
        mc1_chif_ctl_ch3: in     vl_logic_vector(207 downto 0);
        mc1_qif_ctl     : in     vl_logic_vector(143 downto 0);
        pcie_connect    : in     vl_logic_vector(3 downto 0);
        pcie_det_done   : in     vl_logic_vector(3 downto 0);
        pcie_powerdown_ch0: in     vl_logic_vector(1 downto 0);
        pcie_powerdown_ch1: in     vl_logic_vector(1 downto 0);
        pcie_powerdown_ch2: in     vl_logic_vector(1 downto 0);
        pcie_powerdown_ch3: in     vl_logic_vector(1 downto 0);
        pcie_rxpolarity : in     vl_logic_vector(3 downto 0);
        pcie_txcompliance: in     vl_logic_vector(3 downto 0);
        pcie_txdetrx_pr2tlb: in     vl_logic_vector(3 downto 0);
        pcie_txelecidle : in     vl_logic_vector(3 downto 0);
        plol            : in     vl_logic;
        rlol            : in     vl_logic_vector(3 downto 0);
        rlos_hi         : in     vl_logic_vector(3 downto 0);
        rlos_lo         : in     vl_logic_vector(3 downto 0);
        rx_i_clk        : in     vl_logic_vector(3 downto 0);
        sb_rx_d_0       : in     vl_logic_vector(9 downto 0);
        sb_rx_d_1       : in     vl_logic_vector(9 downto 0);
        sb_rx_d_2       : in     vl_logic_vector(9 downto 0);
        sb_rx_d_3       : in     vl_logic_vector(9 downto 0);
        sciaddr         : in     vl_logic_vector(5 downto 0);
        scienaux        : in     vl_logic;
        sciench0        : in     vl_logic;
        sciench1        : in     vl_logic;
        sciench2        : in     vl_logic;
        sciench3        : in     vl_logic;
        scird           : in     vl_logic;
        sciselaux       : in     vl_logic;
        sciselch0       : in     vl_logic;
        sciselch1       : in     vl_logic;
        sciselch2       : in     vl_logic;
        sciselch3       : in     vl_logic;
        sciwdata        : in     vl_logic_vector(7 downto 0);
        sciwstn         : in     vl_logic;
        sd_rx_clk       : in     vl_logic_vector(3 downto 0);
        sd_tx_clk       : in     vl_logic_vector(3 downto 0);
        ser_sts_1_qd_25 : in     vl_logic_vector(7 downto 0);
        ser_sts_2_ch_27_0: in     vl_logic_vector(7 downto 0);
        ser_sts_2_ch_27_1: in     vl_logic_vector(7 downto 0);
        ser_sts_2_ch_27_2: in     vl_logic_vector(7 downto 0);
        ser_sts_2_ch_27_3: in     vl_logic_vector(7 downto 0);
        ser_sts_3_ch_28_0: in     vl_logic_vector(7 downto 0);
        ser_sts_3_ch_28_1: in     vl_logic_vector(7 downto 0);
        ser_sts_3_ch_28_2: in     vl_logic_vector(7 downto 0);
        ser_sts_3_ch_28_3: in     vl_logic_vector(7 downto 0);
        ser_sts_3_qd_27 : in     vl_logic_vector(7 downto 0);
        ser_sts_4_ch_29_0: in     vl_logic_vector(7 downto 0);
        ser_sts_4_ch_29_1: in     vl_logic_vector(7 downto 0);
        ser_sts_4_ch_29_2: in     vl_logic_vector(7 downto 0);
        ser_sts_4_ch_29_3: in     vl_logic_vector(7 downto 0);
        ser_sts_4_qd_28 : in     vl_logic_vector(7 downto 0);
        ser_sts_6_ch_2b_0: in     vl_logic_vector(7 downto 0);
        ser_sts_6_ch_2b_1: in     vl_logic_vector(7 downto 0);
        ser_sts_6_ch_2b_2: in     vl_logic_vector(7 downto 0);
        ser_sts_6_ch_2b_3: in     vl_logic_vector(7 downto 0);
        ser_sts_7_ch_2c_0: in     vl_logic_vector(7 downto 0);
        ser_sts_7_ch_2c_1: in     vl_logic_vector(7 downto 0);
        ser_sts_7_ch_2c_2: in     vl_logic_vector(7 downto 0);
        ser_sts_7_ch_2c_3: in     vl_logic_vector(7 downto 0);
        tck_full        : in     vl_logic;
        tri_ion         : in     vl_logic;
        tx_i_clk        : in     vl_logic_vector(3 downto 0);
        bist_report     : out    vl_logic_vector(15 downto 0);
        cout            : out    vl_logic_vector(19 downto 0);
        ebrd_o_clk      : out    vl_logic_vector(3 downto 0);
        fb_o_clk        : out    vl_logic_vector(3 downto 0);
        ff_rx_d_0       : out    vl_logic_vector(23 downto 0);
        ff_rx_d_1       : out    vl_logic_vector(23 downto 0);
        ff_rx_d_2       : out    vl_logic_vector(23 downto 0);
        ff_rx_d_3       : out    vl_logic_vector(23 downto 0);
        ff_rx_f_clk     : out    vl_logic_vector(3 downto 0);
        ff_rx_h_clk     : out    vl_logic_vector(3 downto 0);
        ff_tx_f_clk     : out    vl_logic_vector(3 downto 0);
        ff_tx_h_clk     : out    vl_logic_vector(3 downto 0);
        fff_pci_det_en  : out    vl_logic_vector(3 downto 0);
        ffr_o_clk       : out    vl_logic_vector(3 downto 0);
        ffs_cc_overrun  : out    vl_logic_vector(3 downto 0);
        ffs_cc_underrun : out    vl_logic_vector(3 downto 0);
        ffs_ls_sync_status: out    vl_logic_vector(3 downto 0);
        ffs_rxfbfifo_error: out    vl_logic_vector(3 downto 0);
        ffs_txfbfifo_error: out    vl_logic_vector(3 downto 0);
        ffs_pcie_phystatus: out    vl_logic_vector(3 downto 0);
        ffs_pcie_rxvalid: out    vl_logic_vector(3 downto 0);
        ffs_skp_added   : out    vl_logic_vector(3 downto 0);
        ffs_skp_deleted : out    vl_logic_vector(3 downto 0);
        fft_o_clk       : out    vl_logic_vector(3 downto 0);
        macro_rst       : out    vl_logic;
        macropdb        : out    vl_logic;
        pcie_beacon_en  : out    vl_logic_vector(3 downto 0);
        pcie_mode       : out    vl_logic_vector(3 downto 0);
        quad_reset_all  : out    vl_logic;
        rrst            : out    vl_logic_vector(3 downto 0);
        rx_o_clk        : out    vl_logic_vector(3 downto 0);
        sb_tx_d_0       : out    vl_logic_vector(9 downto 0);
        sb_tx_d_1       : out    vl_logic_vector(9 downto 0);
        sb_tx_d_2       : out    vl_logic_vector(9 downto 0);
        sb_tx_d_3       : out    vl_logic_vector(9 downto 0);
        sciint          : out    vl_logic;
        scirdata        : out    vl_logic_vector(7 downto 0);
        ser_ctl_1_ch_10_0: out    vl_logic_vector(7 downto 0);
        ser_ctl_1_ch_10_1: out    vl_logic_vector(7 downto 0);
        ser_ctl_1_ch_10_2: out    vl_logic_vector(7 downto 0);
        ser_ctl_1_ch_10_3: out    vl_logic_vector(7 downto 0);
        ser_ctl_1_qd_0a : out    vl_logic_vector(7 downto 0);
        ser_ctl_2_ch_11_0: out    vl_logic_vector(7 downto 0);
        ser_ctl_2_ch_11_1: out    vl_logic_vector(7 downto 0);
        ser_ctl_2_ch_11_2: out    vl_logic_vector(7 downto 0);
        ser_ctl_2_ch_11_3: out    vl_logic_vector(7 downto 0);
        ser_ctl_2_qd_0b : out    vl_logic_vector(7 downto 0);
        ser_ctl_3_ch_12_0: out    vl_logic_vector(7 downto 0);
        ser_ctl_3_ch_12_1: out    vl_logic_vector(7 downto 0);
        ser_ctl_3_ch_12_2: out    vl_logic_vector(7 downto 0);
        ser_ctl_3_ch_12_3: out    vl_logic_vector(7 downto 0);
        ser_ctl_3_qd_0c : out    vl_logic_vector(7 downto 0);
        ser_ctl_4_ch_13_0: out    vl_logic_vector(7 downto 0);
        ser_ctl_4_ch_13_1: out    vl_logic_vector(7 downto 0);
        ser_ctl_4_ch_13_2: out    vl_logic_vector(7 downto 0);
        ser_ctl_4_ch_13_3: out    vl_logic_vector(7 downto 0);
        ser_ctl_4_qd_0d : out    vl_logic_vector(7 downto 0);
        ser_ctl_5_ch_14_0: out    vl_logic_vector(7 downto 0);
        ser_ctl_5_ch_14_1: out    vl_logic_vector(7 downto 0);
        ser_ctl_5_ch_14_2: out    vl_logic_vector(7 downto 0);
        ser_ctl_5_ch_14_3: out    vl_logic_vector(7 downto 0);
        ser_ctl_5_qd_0e : out    vl_logic_vector(7 downto 0);
        ser_ctl_6_ch_15_0: out    vl_logic_vector(7 downto 0);
        ser_ctl_6_ch_15_1: out    vl_logic_vector(7 downto 0);
        ser_ctl_6_ch_15_2: out    vl_logic_vector(7 downto 0);
        ser_ctl_6_ch_15_3: out    vl_logic_vector(7 downto 0);
        ser_ctl_7_ch_16_0: out    vl_logic_vector(7 downto 0);
        ser_ctl_7_ch_16_1: out    vl_logic_vector(7 downto 0);
        ser_ctl_7_ch_16_2: out    vl_logic_vector(7 downto 0);
        ser_ctl_7_ch_16_3: out    vl_logic_vector(7 downto 0);
        ser_ch_rst_0    : out    vl_logic_vector(1 downto 0);
        ser_ch_rst_1    : out    vl_logic_vector(1 downto 0);
        ser_ch_rst_2    : out    vl_logic_vector(1 downto 0);
        ser_ch_rst_3    : out    vl_logic_vector(1 downto 0);
        sync_pulse      : out    vl_logic;
        trst            : out    vl_logic;
        tsd_pcie_det_ct : out    vl_logic_vector(3 downto 0);
        tsd_pcie_ei_en  : out    vl_logic_vector(3 downto 0);
        tx_o_clk        : out    vl_logic_vector(3 downto 0)
    );
end pcs_quad;
