library verilog;
use verilog.vl_types.all;
entity pcs_quad_dp is
    port(
        bus8bit_sel     : in     vl_logic;
        bist_rx_data_sel: in     vl_logic;
        char_mode       : in     vl_logic;
        char_test_data  : in     vl_logic_vector(9 downto 0);
        char_test_mode  : in     vl_logic;
        ebrd_i_clk      : in     vl_logic_vector(3 downto 0);
        fb_i_clk        : in     vl_logic_vector(3 downto 0);
        ff_ebrd_clk     : in     vl_logic_vector(3 downto 0);
        ff_rxi_clk      : in     vl_logic_vector(3 downto 0);
        ff_tx_d_0       : in     vl_logic_vector(23 downto 0);
        ff_tx_d_1       : in     vl_logic_vector(23 downto 0);
        ff_tx_d_2       : in     vl_logic_vector(23 downto 0);
        ff_tx_d_3       : in     vl_logic_vector(23 downto 0);
        ff_txi_clk      : in     vl_logic_vector(3 downto 0);
        ffc_ei_en       : in     vl_logic_vector(3 downto 0);
        ffc_enable_cgalign: in     vl_logic_vector(3 downto 0);
        ffc_fb_loopback : in     vl_logic_vector(3 downto 0);
        ffc_lane_rx_rst : in     vl_logic_vector(3 downto 0);
        ffc_lane_tx_rst : in     vl_logic_vector(3 downto 0);
        ffc_pci_det_en  : in     vl_logic_vector(3 downto 0);
        ffc_pcie_ct     : in     vl_logic_vector(3 downto 0);
        ffc_pfifo_clr   : in     vl_logic_vector(3 downto 0);
        ffc_rxpwdnb     : in     vl_logic_vector(3 downto 0);
        ffc_sb_inv_rx   : in     vl_logic_vector(3 downto 0);
        ffc_sb_pfifo_lp : in     vl_logic_vector(3 downto 0);
        ffc_signal_detect: in     vl_logic_vector(3 downto 0);
        ffc_txpwdnb     : in     vl_logic_vector(3 downto 0);
        ffc_rx_div11_clk: in     vl_logic_vector(3 downto 0);
        ffc_tx_div11_clk: in     vl_logic_vector(3 downto 0);
        ffc_rx_rate_mode: in     vl_logic_vector(3 downto 0);
        ffc_tx_rate_mode: in     vl_logic_vector(3 downto 0);
        ffr_i_clk       : in     vl_logic_vector(3 downto 0);
        fft_i_clk       : in     vl_logic_vector(3 downto 0);
        fmbist_data_0   : in     vl_logic_vector(9 downto 0);
        fmbist_data_1   : in     vl_logic_vector(9 downto 0);
        fmbist_data_2   : in     vl_logic_vector(9 downto 0);
        fmbist_data_3   : in     vl_logic_vector(9 downto 0);
        force_int       : in     vl_logic;
        ffc_ldr_core2tx_en: in     vl_logic_vector(3 downto 0);
        mc1_chif_ctl_ch0: in     vl_logic_vector(207 downto 0);
        mc1_chif_ctl_ch1: in     vl_logic_vector(207 downto 0);
        mc1_chif_ctl_ch2: in     vl_logic_vector(207 downto 0);
        mc1_chif_ctl_ch3: in     vl_logic_vector(207 downto 0);
        pcie_connect    : in     vl_logic_vector(3 downto 0);
        pcie_det_done   : in     vl_logic_vector(3 downto 0);
        pcie_powerdown_ch0: in     vl_logic_vector(1 downto 0);
        pcie_powerdown_ch1: in     vl_logic_vector(1 downto 0);
        pcie_powerdown_ch2: in     vl_logic_vector(1 downto 0);
        pcie_powerdown_ch3: in     vl_logic_vector(1 downto 0);
        pcie_rxpolarity : in     vl_logic_vector(3 downto 0);
        pcie_txcompliance: in     vl_logic_vector(3 downto 0);
        pcie_txdetrx_pr2tlb: in     vl_logic_vector(3 downto 0);
        pcie_txelecidle : in     vl_logic_vector(3 downto 0);
        pcs_ctl_3_qd_02 : in     vl_logic_vector(7 downto 0);
        pcs_ctl_4_qd_03 : in     vl_logic_vector(7 downto 0);
        plol            : in     vl_logic;
        quad_reset_all  : in     vl_logic;
        quad_reset_all_n: in     vl_logic;
        rlol            : in     vl_logic_vector(3 downto 0);
        rlos_hi         : in     vl_logic_vector(3 downto 0);
        rlos_lo         : in     vl_logic_vector(3 downto 0);
        rx_i_clk        : in     vl_logic_vector(3 downto 0);
        sb_rx_d_0       : in     vl_logic_vector(9 downto 0);
        sb_rx_d_1       : in     vl_logic_vector(9 downto 0);
        sb_rx_d_2       : in     vl_logic_vector(9 downto 0);
        sb_rx_d_3       : in     vl_logic_vector(9 downto 0);
        sci_addr10      : in     vl_logic_vector(5 downto 0);
        sci_addr32      : in     vl_logic_vector(5 downto 0);
        sci_ion_dl10    : in     vl_logic;
        sci_ion_dl32    : in     vl_logic;
        sci_rd10        : in     vl_logic;
        sci_rd32        : in     vl_logic;
        sci_resetn10    : in     vl_logic;
        sci_resetn32    : in     vl_logic;
        sci_wdata10     : in     vl_logic_vector(7 downto 0);
        sci_wdata32     : in     vl_logic_vector(7 downto 0);
        sci_wstb10      : in     vl_logic;
        sci_wstb32      : in     vl_logic;
        sciench0_b      : in     vl_logic;
        sciench1_b      : in     vl_logic;
        sciench2_b      : in     vl_logic;
        sciench3_b      : in     vl_logic;
        sciselch0_b     : in     vl_logic;
        sciselch1_b     : in     vl_logic;
        sciselch2_b     : in     vl_logic;
        sciselch3_b     : in     vl_logic;
        sd_rx_clk       : in     vl_logic_vector(3 downto 0);
        sd_tx_clk       : in     vl_logic_vector(3 downto 0);
        ser_sts_2_ch_27_0: in     vl_logic_vector(7 downto 0);
        ser_sts_2_ch_27_1: in     vl_logic_vector(7 downto 0);
        ser_sts_2_ch_27_2: in     vl_logic_vector(7 downto 0);
        ser_sts_2_ch_27_3: in     vl_logic_vector(7 downto 0);
        ser_sts_3_ch_28_0: in     vl_logic_vector(7 downto 0);
        ser_sts_3_ch_28_1: in     vl_logic_vector(7 downto 0);
        ser_sts_3_ch_28_2: in     vl_logic_vector(7 downto 0);
        ser_sts_3_ch_28_3: in     vl_logic_vector(7 downto 0);
        ser_sts_4_ch_29_0: in     vl_logic_vector(7 downto 0);
        ser_sts_4_ch_29_1: in     vl_logic_vector(7 downto 0);
        ser_sts_4_ch_29_2: in     vl_logic_vector(7 downto 0);
        ser_sts_4_ch_29_3: in     vl_logic_vector(7 downto 0);
        ser_sts_6_ch_2b_0: in     vl_logic_vector(7 downto 0);
        ser_sts_6_ch_2b_1: in     vl_logic_vector(7 downto 0);
        ser_sts_6_ch_2b_2: in     vl_logic_vector(7 downto 0);
        ser_sts_6_ch_2b_3: in     vl_logic_vector(7 downto 0);
        ser_sts_7_ch_2c_0: in     vl_logic_vector(7 downto 0);
        ser_sts_7_ch_2c_1: in     vl_logic_vector(7 downto 0);
        ser_sts_7_ch_2c_2: in     vl_logic_vector(7 downto 0);
        ser_sts_7_ch_2c_3: in     vl_logic_vector(7 downto 0);
        test_clk        : in     vl_logic;
        tx_i_clk        : in     vl_logic_vector(3 downto 0);
        xge_mode        : in     vl_logic;
        ebrd_o_clk      : out    vl_logic_vector(3 downto 0);
        fb_o_clk        : out    vl_logic_vector(3 downto 0);
        ff_rx_d_0       : out    vl_logic_vector(23 downto 0);
        ff_rx_d_1       : out    vl_logic_vector(23 downto 0);
        ff_rx_d_2       : out    vl_logic_vector(23 downto 0);
        ff_rx_d_3       : out    vl_logic_vector(23 downto 0);
        ff_rx_f_clk     : out    vl_logic_vector(3 downto 0);
        ff_rx_h_clk     : out    vl_logic_vector(3 downto 0);
        ff_tx_f_clk     : out    vl_logic_vector(3 downto 0);
        ff_tx_h_clk     : out    vl_logic_vector(3 downto 0);
        fff_pci_det_en  : out    vl_logic_vector(3 downto 0);
        ffr_o_clk       : out    vl_logic_vector(3 downto 0);
        ffs_cc_overrun  : out    vl_logic_vector(3 downto 0);
        ffs_cc_underrun : out    vl_logic_vector(3 downto 0);
        ffs_ls_sync_status: out    vl_logic_vector(3 downto 0);
        ffs_rxfbfifo_error: out    vl_logic_vector(3 downto 0);
        ffs_txfbfifo_error: out    vl_logic_vector(3 downto 0);
        fft_o_clk       : out    vl_logic_vector(3 downto 0);
        int_cha_out     : out    vl_logic_vector(3 downto 0);
        pcie_beacon_en  : out    vl_logic_vector(3 downto 0);
        pcie_mode       : out    vl_logic_vector(3 downto 0);
        pcie_phystatus  : out    vl_logic_vector(3 downto 0);
        pcie_rxvalid    : out    vl_logic_vector(3 downto 0);
        skp_added       : out    vl_logic_vector(3 downto 0);
        skp_deleted     : out    vl_logic_vector(3 downto 0);
        rx_ch           : out    vl_logic_vector(3 downto 0);
        rx_o_clk        : out    vl_logic_vector(3 downto 0);
        sb_tx_d_0       : out    vl_logic_vector(9 downto 0);
        sb_tx_d_1       : out    vl_logic_vector(9 downto 0);
        sb_tx_d_2       : out    vl_logic_vector(9 downto 0);
        sb_tx_d_3       : out    vl_logic_vector(9 downto 0);
        sci_int10       : out    vl_logic;
        sci_int32       : out    vl_logic;
        sci_rdata10     : out    vl_logic_vector(7 downto 0);
        sci_rdata32     : out    vl_logic_vector(7 downto 0);
        ser_ctl_1_ch_10_0: out    vl_logic_vector(7 downto 0);
        ser_ctl_1_ch_10_1: out    vl_logic_vector(7 downto 0);
        ser_ctl_1_ch_10_2: out    vl_logic_vector(7 downto 0);
        ser_ctl_1_ch_10_3: out    vl_logic_vector(7 downto 0);
        ser_ctl_2_ch_11_0: out    vl_logic_vector(7 downto 0);
        ser_ctl_2_ch_11_1: out    vl_logic_vector(7 downto 0);
        ser_ctl_2_ch_11_2: out    vl_logic_vector(7 downto 0);
        ser_ctl_2_ch_11_3: out    vl_logic_vector(7 downto 0);
        ser_ctl_3_ch_12_0: out    vl_logic_vector(7 downto 0);
        ser_ctl_3_ch_12_1: out    vl_logic_vector(7 downto 0);
        ser_ctl_3_ch_12_2: out    vl_logic_vector(7 downto 0);
        ser_ctl_3_ch_12_3: out    vl_logic_vector(7 downto 0);
        ser_ctl_4_ch_13_0: out    vl_logic_vector(7 downto 0);
        ser_ctl_4_ch_13_1: out    vl_logic_vector(7 downto 0);
        ser_ctl_4_ch_13_2: out    vl_logic_vector(7 downto 0);
        ser_ctl_4_ch_13_3: out    vl_logic_vector(7 downto 0);
        ser_ctl_5_ch_14_0: out    vl_logic_vector(7 downto 0);
        ser_ctl_5_ch_14_1: out    vl_logic_vector(7 downto 0);
        ser_ctl_5_ch_14_2: out    vl_logic_vector(7 downto 0);
        ser_ctl_5_ch_14_3: out    vl_logic_vector(7 downto 0);
        ser_ctl_6_ch_15_0: out    vl_logic_vector(7 downto 0);
        ser_ctl_6_ch_15_1: out    vl_logic_vector(7 downto 0);
        ser_ctl_6_ch_15_2: out    vl_logic_vector(7 downto 0);
        ser_ctl_6_ch_15_3: out    vl_logic_vector(7 downto 0);
        ser_ctl_7_ch_16_0: out    vl_logic_vector(7 downto 0);
        ser_ctl_7_ch_16_1: out    vl_logic_vector(7 downto 0);
        ser_ctl_7_ch_16_2: out    vl_logic_vector(7 downto 0);
        ser_ctl_7_ch_16_3: out    vl_logic_vector(7 downto 0);
        ser_ch_rst_0    : out    vl_logic_vector(2 downto 0);
        ser_ch_rst_1    : out    vl_logic_vector(2 downto 0);
        ser_ch_rst_2    : out    vl_logic_vector(2 downto 0);
        ser_ch_rst_3    : out    vl_logic_vector(2 downto 0);
        tobist_data_0   : out    vl_logic_vector(9 downto 0);
        tobist_data_1   : out    vl_logic_vector(9 downto 0);
        tobist_data_2   : out    vl_logic_vector(9 downto 0);
        tobist_data_3   : out    vl_logic_vector(9 downto 0);
        tsd_pcie_det_ct : out    vl_logic_vector(3 downto 0);
        tsd_pcie_ei_en  : out    vl_logic_vector(3 downto 0);
        tx_o_clk        : out    vl_logic_vector(3 downto 0)
    );
end pcs_quad_dp;
